module background (
    input [5:0] x_input,
    input [5:0] y_input,
    output [5:0] data
);

logic [11:0] address;
assign address = {y_input, x_input};

always_comb begin
    case(address) 
12'b000000000000: data = 6'b010101;
12'b000000000001: data = 6'b010101;
12'b000000000010: data = 6'b010101;
12'b000000000011: data = 6'b010101;
12'b000000000100: data = 6'b010101;
12'b000000000101: data = 6'b010101;
12'b000000000110: data = 6'b010101;
12'b000000000111: data = 6'b010101;
12'b000000001000: data = 6'b010101;
12'b000000001001: data = 6'b010101;
12'b000000001010: data = 6'b010101;
12'b000000001011: data = 6'b010101;
12'b000000001100: data = 6'b010101;
12'b000000001101: data = 6'b010101;
12'b000000001110: data = 6'b010101;
12'b000000001111: data = 6'b010101;
12'b000000010000: data = 6'b010101;
12'b000000010001: data = 6'b010101;
12'b000000010010: data = 6'b010101;
12'b000000010011: data = 6'b010101;
12'b000000010100: data = 6'b010101;
12'b000000010101: data = 6'b010101;
12'b000000010110: data = 6'b010101;
12'b000000010111: data = 6'b010101;
12'b000000011000: data = 6'b010101;
12'b000000011001: data = 6'b010101;
12'b000000011010: data = 6'b010101;
12'b000000011011: data = 6'b010101;
12'b000000011100: data = 6'b010101;
12'b000000011101: data = 6'b010101;
12'b000000011110: data = 6'b010101;
12'b000000011111: data = 6'b010101;
12'b000000100000: data = 6'b010101;
12'b000000100001: data = 6'b010101;
12'b000000100010: data = 6'b010101;
12'b000000100011: data = 6'b010101;
12'b000000100100: data = 6'b010101;
12'b000000100101: data = 6'b010101;
12'b000000100110: data = 6'b010101;
12'b000000100111: data = 6'b010101;
12'b000000101000: data = 6'b010101;
12'b000000101001: data = 6'b010101;
12'b000000101010: data = 6'b010101;
12'b000000101011: data = 6'b010101;
12'b000000101100: data = 6'b010101;
12'b000000101101: data = 6'b010101;
12'b000000101110: data = 6'b010101;
12'b000000101111: data = 6'b010101;
12'b000000110000: data = 6'b010101;
12'b000000110001: data = 6'b010101;
12'b000000110010: data = 6'b010101;
12'b000000110011: data = 6'b010101;
12'b000000110100: data = 6'b010101;
12'b000000110101: data = 6'b010101;
12'b000000110110: data = 6'b010101;
12'b000000110111: data = 6'b010101;
12'b000000111000: data = 6'b010101;
12'b000000111001: data = 6'b010101;
12'b000000111010: data = 6'b010101;
12'b000000111011: data = 6'b010101;
12'b000000111100: data = 6'b010101;
12'b000000111101: data = 6'b010101;
12'b000000111110: data = 6'b010101;
12'b000000111111: data = 6'b010101;
12'b0000001000000: data = 6'b010101;
12'b0000001000001: data = 6'b010101;
12'b0000001000010: data = 6'b010101;
12'b0000001000011: data = 6'b010101;
12'b0000001000100: data = 6'b010101;
12'b0000001000101: data = 6'b010101;
12'b0000001000110: data = 6'b010101;
12'b0000001000111: data = 6'b010101;
12'b0000001001000: data = 6'b010101;
12'b0000001001001: data = 6'b010101;
12'b0000001001010: data = 6'b010101;
12'b0000001001011: data = 6'b010101;
12'b0000001001100: data = 6'b010101;
12'b0000001001101: data = 6'b010101;
12'b0000001001110: data = 6'b010101;
12'b0000001001111: data = 6'b010101;
12'b0000001010000: data = 6'b010101;
12'b0000001010001: data = 6'b010101;
12'b0000001010010: data = 6'b010101;
12'b0000001010011: data = 6'b010101;
12'b0000001010100: data = 6'b010101;
12'b0000001010101: data = 6'b010101;
12'b0000001010110: data = 6'b010101;
12'b0000001010111: data = 6'b010101;
12'b0000001011000: data = 6'b010101;
12'b0000001011001: data = 6'b010101;
12'b0000001011010: data = 6'b010101;
12'b0000001011011: data = 6'b010101;
12'b0000001011100: data = 6'b010101;
12'b0000001011101: data = 6'b010101;
12'b0000001011110: data = 6'b010101;
12'b0000001011111: data = 6'b010101;
12'b0000001100000: data = 6'b010101;
12'b0000001100001: data = 6'b010101;
12'b0000001100010: data = 6'b010101;
12'b0000001100011: data = 6'b010101;
12'b0000001100100: data = 6'b010101;
12'b0000001100101: data = 6'b010101;
12'b0000001100110: data = 6'b010101;
12'b0000001100111: data = 6'b010101;
12'b0000001101000: data = 6'b010101;
12'b0000001101001: data = 6'b010101;
12'b0000001101010: data = 6'b010101;
12'b0000001101011: data = 6'b010101;
12'b0000001101100: data = 6'b010101;
12'b0000001101101: data = 6'b010101;
12'b0000001101110: data = 6'b010101;
12'b0000001101111: data = 6'b010101;
12'b0000001110000: data = 6'b010101;
12'b0000001110001: data = 6'b010101;
12'b0000001110010: data = 6'b010101;
12'b0000001110011: data = 6'b010101;
12'b0000001110100: data = 6'b010101;
12'b0000001110101: data = 6'b010101;
12'b0000001110110: data = 6'b010101;
12'b0000001110111: data = 6'b010101;
12'b0000001111000: data = 6'b010101;
12'b0000001111001: data = 6'b010101;
12'b0000001111010: data = 6'b010101;
12'b0000001111011: data = 6'b010101;
12'b0000001111100: data = 6'b010101;
12'b0000001111101: data = 6'b010101;
12'b0000001111110: data = 6'b010101;
12'b0000001111111: data = 6'b010101;
12'b00000010000000: data = 6'b010101;
12'b00000010000001: data = 6'b010101;
12'b00000010000010: data = 6'b010101;
12'b00000010000011: data = 6'b010101;
12'b00000010000100: data = 6'b010101;
12'b00000010000101: data = 6'b010101;
12'b00000010000110: data = 6'b010101;
12'b00000010000111: data = 6'b010101;
12'b00000010001000: data = 6'b010101;
12'b00000010001001: data = 6'b010101;
12'b00000010001010: data = 6'b010101;
12'b00000010001011: data = 6'b010101;
12'b00000010001100: data = 6'b010101;
12'b00000010001101: data = 6'b010101;
12'b00000010001110: data = 6'b010101;
12'b00000010001111: data = 6'b010101;
12'b00000010010000: data = 6'b010101;
12'b00000010010001: data = 6'b010101;
12'b00000010010010: data = 6'b010101;
12'b00000010010011: data = 6'b010101;
12'b00000010010100: data = 6'b010101;
12'b00000010010101: data = 6'b010101;
12'b00000010010110: data = 6'b010101;
12'b00000010010111: data = 6'b010101;
12'b00000010011000: data = 6'b010101;
12'b00000010011001: data = 6'b010101;
12'b00000010011010: data = 6'b010101;
12'b00000010011011: data = 6'b010101;
12'b00000010011100: data = 6'b010101;
12'b00000010011101: data = 6'b010101;
12'b00000010011110: data = 6'b010101;
12'b00000010011111: data = 6'b010101;
12'b00000010100000: data = 6'b010101;
12'b00000010100001: data = 6'b010101;
12'b00000010100010: data = 6'b010101;
12'b00000010100011: data = 6'b010101;
12'b00000010100100: data = 6'b010101;
12'b00000010100101: data = 6'b010101;
12'b00000010100110: data = 6'b010101;
12'b00000010100111: data = 6'b010101;
12'b00000010101000: data = 6'b010101;
12'b00000010101001: data = 6'b010101;
12'b00000010101010: data = 6'b010101;
12'b000001000000: data = 6'b010101;
12'b000001000001: data = 6'b010101;
12'b000001000010: data = 6'b010101;
12'b000001000011: data = 6'b010101;
12'b000001000100: data = 6'b010101;
12'b000001000101: data = 6'b010101;
12'b000001000110: data = 6'b010101;
12'b000001000111: data = 6'b010101;
12'b000001001000: data = 6'b010101;
12'b000001001001: data = 6'b010101;
12'b000001001010: data = 6'b010101;
12'b000001001011: data = 6'b010101;
12'b000001001100: data = 6'b010101;
12'b000001001101: data = 6'b010101;
12'b000001001110: data = 6'b010101;
12'b000001001111: data = 6'b010101;
12'b000001010000: data = 6'b010101;
12'b000001010001: data = 6'b010101;
12'b000001010010: data = 6'b010101;
12'b000001010011: data = 6'b010101;
12'b000001010100: data = 6'b010101;
12'b000001010101: data = 6'b010101;
12'b000001010110: data = 6'b010101;
12'b000001010111: data = 6'b010101;
12'b000001011000: data = 6'b010101;
12'b000001011001: data = 6'b010101;
12'b000001011010: data = 6'b010101;
12'b000001011011: data = 6'b010101;
12'b000001011100: data = 6'b010101;
12'b000001011101: data = 6'b010101;
12'b000001011110: data = 6'b010101;
12'b000001011111: data = 6'b010101;
12'b000001100000: data = 6'b010101;
12'b000001100001: data = 6'b010101;
12'b000001100010: data = 6'b010101;
12'b000001100011: data = 6'b010101;
12'b000001100100: data = 6'b010101;
12'b000001100101: data = 6'b010101;
12'b000001100110: data = 6'b010101;
12'b000001100111: data = 6'b010101;
12'b000001101000: data = 6'b010101;
12'b000001101001: data = 6'b010101;
12'b000001101010: data = 6'b010101;
12'b000001101011: data = 6'b010101;
12'b000001101100: data = 6'b010101;
12'b000001101101: data = 6'b010101;
12'b000001101110: data = 6'b010101;
12'b000001101111: data = 6'b010101;
12'b000001110000: data = 6'b010101;
12'b000001110001: data = 6'b010101;
12'b000001110010: data = 6'b010101;
12'b000001110011: data = 6'b010101;
12'b000001110100: data = 6'b010101;
12'b000001110101: data = 6'b010101;
12'b000001110110: data = 6'b010101;
12'b000001110111: data = 6'b010101;
12'b000001111000: data = 6'b010101;
12'b000001111001: data = 6'b010101;
12'b000001111010: data = 6'b010101;
12'b000001111011: data = 6'b010101;
12'b000001111100: data = 6'b010101;
12'b000001111101: data = 6'b010101;
12'b000001111110: data = 6'b010101;
12'b000001111111: data = 6'b010101;
12'b0000011000000: data = 6'b010101;
12'b0000011000001: data = 6'b010101;
12'b0000011000010: data = 6'b010101;
12'b0000011000011: data = 6'b010101;
12'b0000011000100: data = 6'b010101;
12'b0000011000101: data = 6'b010101;
12'b0000011000110: data = 6'b010101;
12'b0000011000111: data = 6'b010101;
12'b0000011001000: data = 6'b010101;
12'b0000011001001: data = 6'b010101;
12'b0000011001010: data = 6'b010101;
12'b0000011001011: data = 6'b010101;
12'b0000011001100: data = 6'b010101;
12'b0000011001101: data = 6'b010101;
12'b0000011001110: data = 6'b010101;
12'b0000011001111: data = 6'b010101;
12'b0000011010000: data = 6'b010101;
12'b0000011010001: data = 6'b010101;
12'b0000011010010: data = 6'b010101;
12'b0000011010011: data = 6'b010101;
12'b0000011010100: data = 6'b010101;
12'b0000011010101: data = 6'b010101;
12'b0000011010110: data = 6'b010101;
12'b0000011010111: data = 6'b010101;
12'b0000011011000: data = 6'b010101;
12'b0000011011001: data = 6'b010101;
12'b0000011011010: data = 6'b010101;
12'b0000011011011: data = 6'b010101;
12'b0000011011100: data = 6'b010101;
12'b0000011011101: data = 6'b010101;
12'b0000011011110: data = 6'b010101;
12'b0000011011111: data = 6'b010101;
12'b0000011100000: data = 6'b010101;
12'b0000011100001: data = 6'b010101;
12'b0000011100010: data = 6'b010101;
12'b0000011100011: data = 6'b010101;
12'b0000011100100: data = 6'b010101;
12'b0000011100101: data = 6'b010101;
12'b0000011100110: data = 6'b010101;
12'b0000011100111: data = 6'b010101;
12'b0000011101000: data = 6'b010101;
12'b0000011101001: data = 6'b010101;
12'b0000011101010: data = 6'b010101;
12'b0000011101011: data = 6'b010101;
12'b0000011101100: data = 6'b010101;
12'b0000011101101: data = 6'b010101;
12'b0000011101110: data = 6'b010101;
12'b0000011101111: data = 6'b010101;
12'b0000011110000: data = 6'b010101;
12'b0000011110001: data = 6'b010101;
12'b0000011110010: data = 6'b010101;
12'b0000011110011: data = 6'b010101;
12'b0000011110100: data = 6'b010101;
12'b0000011110101: data = 6'b010101;
12'b0000011110110: data = 6'b010101;
12'b0000011110111: data = 6'b010101;
12'b0000011111000: data = 6'b010101;
12'b0000011111001: data = 6'b010101;
12'b0000011111010: data = 6'b010101;
12'b0000011111011: data = 6'b010101;
12'b0000011111100: data = 6'b010101;
12'b0000011111101: data = 6'b010101;
12'b0000011111110: data = 6'b010101;
12'b0000011111111: data = 6'b010101;
12'b00000110000000: data = 6'b010101;
12'b00000110000001: data = 6'b010101;
12'b00000110000010: data = 6'b010101;
12'b00000110000011: data = 6'b010101;
12'b00000110000100: data = 6'b010101;
12'b00000110000101: data = 6'b010101;
12'b00000110000110: data = 6'b010101;
12'b00000110000111: data = 6'b010101;
12'b00000110001000: data = 6'b010101;
12'b00000110001001: data = 6'b010101;
12'b00000110001010: data = 6'b010101;
12'b00000110001011: data = 6'b010101;
12'b00000110001100: data = 6'b010101;
12'b00000110001101: data = 6'b010101;
12'b00000110001110: data = 6'b010101;
12'b00000110001111: data = 6'b010101;
12'b00000110010000: data = 6'b010101;
12'b00000110010001: data = 6'b010101;
12'b00000110010010: data = 6'b010101;
12'b00000110010011: data = 6'b010101;
12'b00000110010100: data = 6'b010101;
12'b00000110010101: data = 6'b010101;
12'b00000110010110: data = 6'b010101;
12'b00000110010111: data = 6'b010101;
12'b00000110011000: data = 6'b010101;
12'b00000110011001: data = 6'b010101;
12'b00000110011010: data = 6'b010101;
12'b00000110011011: data = 6'b010101;
12'b00000110011100: data = 6'b010101;
12'b00000110011101: data = 6'b010101;
12'b00000110011110: data = 6'b010101;
12'b00000110011111: data = 6'b010101;
12'b00000110100000: data = 6'b010101;
12'b00000110100001: data = 6'b010101;
12'b00000110100010: data = 6'b010101;
12'b00000110100011: data = 6'b010101;
12'b00000110100100: data = 6'b010101;
12'b00000110100101: data = 6'b010101;
12'b00000110100110: data = 6'b010101;
12'b00000110100111: data = 6'b010101;
12'b00000110101000: data = 6'b010101;
12'b00000110101001: data = 6'b010101;
12'b00000110101010: data = 6'b010101;
12'b000010000000: data = 6'b010101;
12'b000010000001: data = 6'b010101;
12'b000010000010: data = 6'b010101;
12'b000010000011: data = 6'b010101;
12'b000010000100: data = 6'b010101;
12'b000010000101: data = 6'b010101;
12'b000010000110: data = 6'b010101;
12'b000010000111: data = 6'b010101;
12'b000010001000: data = 6'b010101;
12'b000010001001: data = 6'b010101;
12'b000010001010: data = 6'b010101;
12'b000010001011: data = 6'b010101;
12'b000010001100: data = 6'b010101;
12'b000010001101: data = 6'b010101;
12'b000010001110: data = 6'b010101;
12'b000010001111: data = 6'b010101;
12'b000010010000: data = 6'b010101;
12'b000010010001: data = 6'b010101;
12'b000010010010: data = 6'b010101;
12'b000010010011: data = 6'b010101;
12'b000010010100: data = 6'b010101;
12'b000010010101: data = 6'b010101;
12'b000010010110: data = 6'b010101;
12'b000010010111: data = 6'b010101;
12'b000010011000: data = 6'b010101;
12'b000010011001: data = 6'b010101;
12'b000010011010: data = 6'b010101;
12'b000010011011: data = 6'b010101;
12'b000010011100: data = 6'b010101;
12'b000010011101: data = 6'b010101;
12'b000010011110: data = 6'b010101;
12'b000010011111: data = 6'b010101;
12'b000010100000: data = 6'b010101;
12'b000010100001: data = 6'b010101;
12'b000010100010: data = 6'b010101;
12'b000010100011: data = 6'b010101;
12'b000010100100: data = 6'b010101;
12'b000010100101: data = 6'b010101;
12'b000010100110: data = 6'b010101;
12'b000010100111: data = 6'b010101;
12'b000010101000: data = 6'b010101;
12'b000010101001: data = 6'b010101;
12'b000010101010: data = 6'b010101;
12'b000010101011: data = 6'b010101;
12'b000010101100: data = 6'b010101;
12'b000010101101: data = 6'b010101;
12'b000010101110: data = 6'b010101;
12'b000010101111: data = 6'b010101;
12'b000010110000: data = 6'b010101;
12'b000010110001: data = 6'b010101;
12'b000010110010: data = 6'b010101;
12'b000010110011: data = 6'b010101;
12'b000010110100: data = 6'b010101;
12'b000010110101: data = 6'b010101;
12'b000010110110: data = 6'b010101;
12'b000010110111: data = 6'b010101;
12'b000010111000: data = 6'b010101;
12'b000010111001: data = 6'b010101;
12'b000010111010: data = 6'b010101;
12'b000010111011: data = 6'b010101;
12'b000010111100: data = 6'b010101;
12'b000010111101: data = 6'b010101;
12'b000010111110: data = 6'b010101;
12'b000010111111: data = 6'b010101;
12'b0000101000000: data = 6'b010101;
12'b0000101000001: data = 6'b010101;
12'b0000101000010: data = 6'b010101;
12'b0000101000011: data = 6'b010101;
12'b0000101000100: data = 6'b010101;
12'b0000101000101: data = 6'b010101;
12'b0000101000110: data = 6'b010101;
12'b0000101000111: data = 6'b010101;
12'b0000101001000: data = 6'b010101;
12'b0000101001001: data = 6'b010101;
12'b0000101001010: data = 6'b010101;
12'b0000101001011: data = 6'b010101;
12'b0000101001100: data = 6'b010101;
12'b0000101001101: data = 6'b010101;
12'b0000101001110: data = 6'b010101;
12'b0000101001111: data = 6'b010101;
12'b0000101010000: data = 6'b010101;
12'b0000101010001: data = 6'b010101;
12'b0000101010010: data = 6'b010101;
12'b0000101010011: data = 6'b010101;
12'b0000101010100: data = 6'b010101;
12'b0000101010101: data = 6'b010101;
12'b0000101010110: data = 6'b010101;
12'b0000101010111: data = 6'b010101;
12'b0000101011000: data = 6'b010101;
12'b0000101011001: data = 6'b010101;
12'b0000101011010: data = 6'b010101;
12'b0000101011011: data = 6'b010101;
12'b0000101011100: data = 6'b010101;
12'b0000101011101: data = 6'b010101;
12'b0000101011110: data = 6'b010101;
12'b0000101011111: data = 6'b010101;
12'b0000101100000: data = 6'b010101;
12'b0000101100001: data = 6'b010101;
12'b0000101100010: data = 6'b010101;
12'b0000101100011: data = 6'b010101;
12'b0000101100100: data = 6'b010101;
12'b0000101100101: data = 6'b010101;
12'b0000101100110: data = 6'b010101;
12'b0000101100111: data = 6'b010101;
12'b0000101101000: data = 6'b010101;
12'b0000101101001: data = 6'b010101;
12'b0000101101010: data = 6'b010101;
12'b0000101101011: data = 6'b010101;
12'b0000101101100: data = 6'b010101;
12'b0000101101101: data = 6'b010101;
12'b0000101101110: data = 6'b010101;
12'b0000101101111: data = 6'b010101;
12'b0000101110000: data = 6'b010101;
12'b0000101110001: data = 6'b010101;
12'b0000101110010: data = 6'b010101;
12'b0000101110011: data = 6'b010101;
12'b0000101110100: data = 6'b010101;
12'b0000101110101: data = 6'b010101;
12'b0000101110110: data = 6'b010101;
12'b0000101110111: data = 6'b010101;
12'b0000101111000: data = 6'b010101;
12'b0000101111001: data = 6'b010101;
12'b0000101111010: data = 6'b010101;
12'b0000101111011: data = 6'b010101;
12'b0000101111100: data = 6'b010101;
12'b0000101111101: data = 6'b010101;
12'b0000101111110: data = 6'b010101;
12'b0000101111111: data = 6'b010101;
12'b00001010000000: data = 6'b010101;
12'b00001010000001: data = 6'b010101;
12'b00001010000010: data = 6'b010101;
12'b00001010000011: data = 6'b010101;
12'b00001010000100: data = 6'b010101;
12'b00001010000101: data = 6'b010101;
12'b00001010000110: data = 6'b010101;
12'b00001010000111: data = 6'b010101;
12'b00001010001000: data = 6'b010101;
12'b00001010001001: data = 6'b010101;
12'b00001010001010: data = 6'b010101;
12'b00001010001011: data = 6'b101010;
12'b00001010001100: data = 6'b101010;
12'b00001010001101: data = 6'b101010;
12'b00001010001110: data = 6'b010101;
12'b00001010001111: data = 6'b010101;
12'b00001010010000: data = 6'b010101;
12'b00001010010001: data = 6'b010101;
12'b00001010010010: data = 6'b010101;
12'b00001010010011: data = 6'b010101;
12'b00001010010100: data = 6'b010101;
12'b00001010010101: data = 6'b010101;
12'b00001010010110: data = 6'b010101;
12'b00001010010111: data = 6'b010101;
12'b00001010011000: data = 6'b010101;
12'b00001010011001: data = 6'b010101;
12'b00001010011010: data = 6'b010101;
12'b00001010011011: data = 6'b010101;
12'b00001010011100: data = 6'b010101;
12'b00001010011101: data = 6'b010101;
12'b00001010011110: data = 6'b010101;
12'b00001010011111: data = 6'b010101;
12'b00001010100000: data = 6'b010101;
12'b00001010100001: data = 6'b010101;
12'b00001010100010: data = 6'b010101;
12'b00001010100011: data = 6'b010101;
12'b00001010100100: data = 6'b010101;
12'b00001010100101: data = 6'b010101;
12'b00001010100110: data = 6'b010101;
12'b00001010100111: data = 6'b010101;
12'b00001010101000: data = 6'b010101;
12'b00001010101001: data = 6'b010101;
12'b00001010101010: data = 6'b010101;
12'b000011000000: data = 6'b010101;
12'b000011000001: data = 6'b010101;
12'b000011000010: data = 6'b010101;
12'b000011000011: data = 6'b010101;
12'b000011000100: data = 6'b010101;
12'b000011000101: data = 6'b010101;
12'b000011000110: data = 6'b010101;
12'b000011000111: data = 6'b010101;
12'b000011001000: data = 6'b010101;
12'b000011001001: data = 6'b010101;
12'b000011001010: data = 6'b010101;
12'b000011001011: data = 6'b010101;
12'b000011001100: data = 6'b010101;
12'b000011001101: data = 6'b010101;
12'b000011001110: data = 6'b010101;
12'b000011001111: data = 6'b010101;
12'b000011010000: data = 6'b010101;
12'b000011010001: data = 6'b010101;
12'b000011010010: data = 6'b010101;
12'b000011010011: data = 6'b010101;
12'b000011010100: data = 6'b010101;
12'b000011010101: data = 6'b010101;
12'b000011010110: data = 6'b010101;
12'b000011010111: data = 6'b010101;
12'b000011011000: data = 6'b010101;
12'b000011011001: data = 6'b010101;
12'b000011011010: data = 6'b010101;
12'b000011011011: data = 6'b010101;
12'b000011011100: data = 6'b010101;
12'b000011011101: data = 6'b010101;
12'b000011011110: data = 6'b010101;
12'b000011011111: data = 6'b010101;
12'b000011100000: data = 6'b010101;
12'b000011100001: data = 6'b010101;
12'b000011100010: data = 6'b010101;
12'b000011100011: data = 6'b010101;
12'b000011100100: data = 6'b010101;
12'b000011100101: data = 6'b010101;
12'b000011100110: data = 6'b010101;
12'b000011100111: data = 6'b010101;
12'b000011101000: data = 6'b010101;
12'b000011101001: data = 6'b010101;
12'b000011101010: data = 6'b010101;
12'b000011101011: data = 6'b010101;
12'b000011101100: data = 6'b010101;
12'b000011101101: data = 6'b010101;
12'b000011101110: data = 6'b010101;
12'b000011101111: data = 6'b010101;
12'b000011110000: data = 6'b010101;
12'b000011110001: data = 6'b010101;
12'b000011110010: data = 6'b010101;
12'b000011110011: data = 6'b010101;
12'b000011110100: data = 6'b010101;
12'b000011110101: data = 6'b010101;
12'b000011110110: data = 6'b010101;
12'b000011110111: data = 6'b010101;
12'b000011111000: data = 6'b010101;
12'b000011111001: data = 6'b010101;
12'b000011111010: data = 6'b010101;
12'b000011111011: data = 6'b010101;
12'b000011111100: data = 6'b010101;
12'b000011111101: data = 6'b010101;
12'b000011111110: data = 6'b010101;
12'b000011111111: data = 6'b010101;
12'b0000111000000: data = 6'b010101;
12'b0000111000001: data = 6'b010101;
12'b0000111000010: data = 6'b010101;
12'b0000111000011: data = 6'b010101;
12'b0000111000100: data = 6'b010101;
12'b0000111000101: data = 6'b010101;
12'b0000111000110: data = 6'b010101;
12'b0000111000111: data = 6'b010101;
12'b0000111001000: data = 6'b010101;
12'b0000111001001: data = 6'b010101;
12'b0000111001010: data = 6'b010101;
12'b0000111001011: data = 6'b010101;
12'b0000111001100: data = 6'b010101;
12'b0000111001101: data = 6'b010101;
12'b0000111001110: data = 6'b010101;
12'b0000111001111: data = 6'b010101;
12'b0000111010000: data = 6'b010101;
12'b0000111010001: data = 6'b010101;
12'b0000111010010: data = 6'b010101;
12'b0000111010011: data = 6'b010101;
12'b0000111010100: data = 6'b010101;
12'b0000111010101: data = 6'b010101;
12'b0000111010110: data = 6'b010101;
12'b0000111010111: data = 6'b010101;
12'b0000111011000: data = 6'b010101;
12'b0000111011001: data = 6'b010101;
12'b0000111011010: data = 6'b010101;
12'b0000111011011: data = 6'b010101;
12'b0000111011100: data = 6'b010101;
12'b0000111011101: data = 6'b010101;
12'b0000111011110: data = 6'b010101;
12'b0000111011111: data = 6'b010101;
12'b0000111100000: data = 6'b010101;
12'b0000111100001: data = 6'b010101;
12'b0000111100010: data = 6'b010101;
12'b0000111100011: data = 6'b010101;
12'b0000111100100: data = 6'b010101;
12'b0000111100101: data = 6'b010101;
12'b0000111100110: data = 6'b010101;
12'b0000111100111: data = 6'b010101;
12'b0000111101000: data = 6'b010101;
12'b0000111101001: data = 6'b010101;
12'b0000111101010: data = 6'b010101;
12'b0000111101011: data = 6'b010101;
12'b0000111101100: data = 6'b010101;
12'b0000111101101: data = 6'b010101;
12'b0000111101110: data = 6'b010101;
12'b0000111101111: data = 6'b010101;
12'b0000111110000: data = 6'b010101;
12'b0000111110001: data = 6'b010101;
12'b0000111110010: data = 6'b010101;
12'b0000111110011: data = 6'b010101;
12'b0000111110100: data = 6'b010101;
12'b0000111110101: data = 6'b010101;
12'b0000111110110: data = 6'b010101;
12'b0000111110111: data = 6'b010101;
12'b0000111111000: data = 6'b010101;
12'b0000111111001: data = 6'b010101;
12'b0000111111010: data = 6'b010101;
12'b0000111111011: data = 6'b010101;
12'b0000111111100: data = 6'b010101;
12'b0000111111101: data = 6'b010101;
12'b0000111111110: data = 6'b010101;
12'b0000111111111: data = 6'b010101;
12'b00001110000000: data = 6'b010101;
12'b00001110000001: data = 6'b010101;
12'b00001110000010: data = 6'b010101;
12'b00001110000011: data = 6'b010101;
12'b00001110000100: data = 6'b010101;
12'b00001110000101: data = 6'b010101;
12'b00001110000110: data = 6'b010101;
12'b00001110000111: data = 6'b010101;
12'b00001110001000: data = 6'b010101;
12'b00001110001001: data = 6'b010101;
12'b00001110001010: data = 6'b010101;
12'b00001110001011: data = 6'b101010;
12'b00001110001100: data = 6'b101010;
12'b00001110001101: data = 6'b101010;
12'b00001110001110: data = 6'b010101;
12'b00001110001111: data = 6'b010101;
12'b00001110010000: data = 6'b010101;
12'b00001110010001: data = 6'b010101;
12'b00001110010010: data = 6'b010101;
12'b00001110010011: data = 6'b010101;
12'b00001110010100: data = 6'b010101;
12'b00001110010101: data = 6'b010101;
12'b00001110010110: data = 6'b010101;
12'b00001110010111: data = 6'b010101;
12'b00001110011000: data = 6'b010101;
12'b00001110011001: data = 6'b010101;
12'b00001110011010: data = 6'b010101;
12'b00001110011011: data = 6'b010101;
12'b00001110011100: data = 6'b010101;
12'b00001110011101: data = 6'b010101;
12'b00001110011110: data = 6'b010101;
12'b00001110011111: data = 6'b010101;
12'b00001110100000: data = 6'b010101;
12'b00001110100001: data = 6'b010101;
12'b00001110100010: data = 6'b010101;
12'b00001110100011: data = 6'b010101;
12'b00001110100100: data = 6'b010101;
12'b00001110100101: data = 6'b010101;
12'b00001110100110: data = 6'b010101;
12'b00001110100111: data = 6'b010101;
12'b00001110101000: data = 6'b010101;
12'b00001110101001: data = 6'b010101;
12'b00001110101010: data = 6'b010101;
12'b000100000000: data = 6'b010101;
12'b000100000001: data = 6'b010101;
12'b000100000010: data = 6'b010101;
12'b000100000011: data = 6'b010101;
12'b000100000100: data = 6'b010101;
12'b000100000101: data = 6'b010101;
12'b000100000110: data = 6'b010101;
12'b000100000111: data = 6'b010101;
12'b000100001000: data = 6'b010101;
12'b000100001001: data = 6'b010101;
12'b000100001010: data = 6'b010101;
12'b000100001011: data = 6'b010101;
12'b000100001100: data = 6'b010101;
12'b000100001101: data = 6'b010101;
12'b000100001110: data = 6'b010101;
12'b000100001111: data = 6'b010101;
12'b000100010000: data = 6'b010101;
12'b000100010001: data = 6'b010101;
12'b000100010010: data = 6'b010101;
12'b000100010011: data = 6'b010101;
12'b000100010100: data = 6'b010101;
12'b000100010101: data = 6'b010101;
12'b000100010110: data = 6'b010101;
12'b000100010111: data = 6'b010101;
12'b000100011000: data = 6'b010101;
12'b000100011001: data = 6'b010101;
12'b000100011010: data = 6'b010101;
12'b000100011011: data = 6'b010101;
12'b000100011100: data = 6'b010101;
12'b000100011101: data = 6'b010101;
12'b000100011110: data = 6'b010101;
12'b000100011111: data = 6'b010101;
12'b000100100000: data = 6'b010101;
12'b000100100001: data = 6'b010101;
12'b000100100010: data = 6'b010101;
12'b000100100011: data = 6'b010101;
12'b000100100100: data = 6'b010101;
12'b000100100101: data = 6'b010101;
12'b000100100110: data = 6'b010101;
12'b000100100111: data = 6'b010101;
12'b000100101000: data = 6'b010101;
12'b000100101001: data = 6'b010101;
12'b000100101010: data = 6'b010101;
12'b000100101011: data = 6'b010101;
12'b000100101100: data = 6'b010101;
12'b000100101101: data = 6'b010101;
12'b000100101110: data = 6'b010101;
12'b000100101111: data = 6'b010101;
12'b000100110000: data = 6'b010101;
12'b000100110001: data = 6'b010101;
12'b000100110010: data = 6'b010101;
12'b000100110011: data = 6'b010101;
12'b000100110100: data = 6'b010101;
12'b000100110101: data = 6'b010101;
12'b000100110110: data = 6'b010101;
12'b000100110111: data = 6'b010101;
12'b000100111000: data = 6'b010101;
12'b000100111001: data = 6'b010101;
12'b000100111010: data = 6'b010101;
12'b000100111011: data = 6'b010101;
12'b000100111100: data = 6'b010101;
12'b000100111101: data = 6'b010101;
12'b000100111110: data = 6'b010101;
12'b000100111111: data = 6'b010101;
12'b0001001000000: data = 6'b010101;
12'b0001001000001: data = 6'b010101;
12'b0001001000010: data = 6'b010101;
12'b0001001000011: data = 6'b010101;
12'b0001001000100: data = 6'b010101;
12'b0001001000101: data = 6'b010101;
12'b0001001000110: data = 6'b010101;
12'b0001001000111: data = 6'b010101;
12'b0001001001000: data = 6'b010101;
12'b0001001001001: data = 6'b010101;
12'b0001001001010: data = 6'b010101;
12'b0001001001011: data = 6'b010101;
12'b0001001001100: data = 6'b010101;
12'b0001001001101: data = 6'b010101;
12'b0001001001110: data = 6'b010101;
12'b0001001001111: data = 6'b010101;
12'b0001001010000: data = 6'b010101;
12'b0001001010001: data = 6'b010101;
12'b0001001010010: data = 6'b010101;
12'b0001001010011: data = 6'b010101;
12'b0001001010100: data = 6'b010101;
12'b0001001010101: data = 6'b010101;
12'b0001001010110: data = 6'b010101;
12'b0001001010111: data = 6'b010101;
12'b0001001011000: data = 6'b010101;
12'b0001001011001: data = 6'b010101;
12'b0001001011010: data = 6'b010101;
12'b0001001011011: data = 6'b010101;
12'b0001001011100: data = 6'b010101;
12'b0001001011101: data = 6'b010101;
12'b0001001011110: data = 6'b010101;
12'b0001001011111: data = 6'b010101;
12'b0001001100000: data = 6'b010101;
12'b0001001100001: data = 6'b010101;
12'b0001001100010: data = 6'b010101;
12'b0001001100011: data = 6'b010101;
12'b0001001100100: data = 6'b010101;
12'b0001001100101: data = 6'b010101;
12'b0001001100110: data = 6'b010101;
12'b0001001100111: data = 6'b010101;
12'b0001001101000: data = 6'b010101;
12'b0001001101001: data = 6'b010101;
12'b0001001101010: data = 6'b010101;
12'b0001001101011: data = 6'b010101;
12'b0001001101100: data = 6'b010101;
12'b0001001101101: data = 6'b010101;
12'b0001001101110: data = 6'b010101;
12'b0001001101111: data = 6'b010101;
12'b0001001110000: data = 6'b010101;
12'b0001001110001: data = 6'b010101;
12'b0001001110010: data = 6'b010101;
12'b0001001110011: data = 6'b010101;
12'b0001001110100: data = 6'b010101;
12'b0001001110101: data = 6'b010101;
12'b0001001110110: data = 6'b010101;
12'b0001001110111: data = 6'b010101;
12'b0001001111000: data = 6'b010101;
12'b0001001111001: data = 6'b010101;
12'b0001001111010: data = 6'b010101;
12'b0001001111011: data = 6'b010101;
12'b0001001111100: data = 6'b010101;
12'b0001001111101: data = 6'b010101;
12'b0001001111110: data = 6'b010101;
12'b0001001111111: data = 6'b010101;
12'b00010010000000: data = 6'b010101;
12'b00010010000001: data = 6'b010101;
12'b00010010000010: data = 6'b010101;
12'b00010010000011: data = 6'b010101;
12'b00010010000100: data = 6'b010101;
12'b00010010000101: data = 6'b010101;
12'b00010010000110: data = 6'b010101;
12'b00010010000111: data = 6'b010101;
12'b00010010001000: data = 6'b010101;
12'b00010010001001: data = 6'b010101;
12'b00010010001010: data = 6'b010101;
12'b00010010001011: data = 6'b010101;
12'b00010010001100: data = 6'b000000;
12'b00010010001101: data = 6'b000000;
12'b00010010001110: data = 6'b010101;
12'b00010010001111: data = 6'b010101;
12'b00010010010000: data = 6'b010101;
12'b00010010010001: data = 6'b010101;
12'b00010010010010: data = 6'b010101;
12'b00010010010011: data = 6'b010101;
12'b00010010010100: data = 6'b010101;
12'b00010010010101: data = 6'b010101;
12'b00010010010110: data = 6'b010101;
12'b00010010010111: data = 6'b010101;
12'b00010010011000: data = 6'b010101;
12'b00010010011001: data = 6'b010101;
12'b00010010011010: data = 6'b010101;
12'b00010010011011: data = 6'b010101;
12'b00010010011100: data = 6'b010101;
12'b00010010011101: data = 6'b010101;
12'b00010010011110: data = 6'b010101;
12'b00010010011111: data = 6'b010101;
12'b00010010100000: data = 6'b010101;
12'b00010010100001: data = 6'b010101;
12'b00010010100010: data = 6'b010101;
12'b00010010100011: data = 6'b010101;
12'b00010010100100: data = 6'b010101;
12'b00010010100101: data = 6'b010101;
12'b00010010100110: data = 6'b010101;
12'b00010010100111: data = 6'b010101;
12'b00010010101000: data = 6'b010101;
12'b00010010101001: data = 6'b010101;
12'b00010010101010: data = 6'b010101;
12'b000101000000: data = 6'b010101;
12'b000101000001: data = 6'b010101;
12'b000101000010: data = 6'b010101;
12'b000101000011: data = 6'b010101;
12'b000101000100: data = 6'b010101;
12'b000101000101: data = 6'b010101;
12'b000101000110: data = 6'b010101;
12'b000101000111: data = 6'b010101;
12'b000101001000: data = 6'b010101;
12'b000101001001: data = 6'b010101;
12'b000101001010: data = 6'b010101;
12'b000101001011: data = 6'b010101;
12'b000101001100: data = 6'b010101;
12'b000101001101: data = 6'b010101;
12'b000101001110: data = 6'b010101;
12'b000101001111: data = 6'b010101;
12'b000101010000: data = 6'b010101;
12'b000101010001: data = 6'b010101;
12'b000101010010: data = 6'b010101;
12'b000101010011: data = 6'b010101;
12'b000101010100: data = 6'b010101;
12'b000101010101: data = 6'b010101;
12'b000101010110: data = 6'b010101;
12'b000101010111: data = 6'b010101;
12'b000101011000: data = 6'b010101;
12'b000101011001: data = 6'b010101;
12'b000101011010: data = 6'b101010;
12'b000101011011: data = 6'b101010;
12'b000101011100: data = 6'b101010;
12'b000101011101: data = 6'b101010;
12'b000101011110: data = 6'b101010;
12'b000101011111: data = 6'b101010;
12'b000101100000: data = 6'b101010;
12'b000101100001: data = 6'b101010;
12'b000101100010: data = 6'b101010;
12'b000101100011: data = 6'b101010;
12'b000101100100: data = 6'b101010;
12'b000101100101: data = 6'b010101;
12'b000101100110: data = 6'b010101;
12'b000101100111: data = 6'b010101;
12'b000101101000: data = 6'b010101;
12'b000101101001: data = 6'b010101;
12'b000101101010: data = 6'b010101;
12'b000101101011: data = 6'b010101;
12'b000101101100: data = 6'b010101;
12'b000101101101: data = 6'b010101;
12'b000101101110: data = 6'b010101;
12'b000101101111: data = 6'b010101;
12'b000101110000: data = 6'b010101;
12'b000101110001: data = 6'b010101;
12'b000101110010: data = 6'b010101;
12'b000101110011: data = 6'b010101;
12'b000101110100: data = 6'b010101;
12'b000101110101: data = 6'b010101;
12'b000101110110: data = 6'b010101;
12'b000101110111: data = 6'b010101;
12'b000101111000: data = 6'b010101;
12'b000101111001: data = 6'b010101;
12'b000101111010: data = 6'b010101;
12'b000101111011: data = 6'b010101;
12'b000101111100: data = 6'b010101;
12'b000101111101: data = 6'b010101;
12'b000101111110: data = 6'b010101;
12'b000101111111: data = 6'b010101;
12'b0001011000000: data = 6'b010101;
12'b0001011000001: data = 6'b010101;
12'b0001011000010: data = 6'b010101;
12'b0001011000011: data = 6'b010101;
12'b0001011000100: data = 6'b010101;
12'b0001011000101: data = 6'b010101;
12'b0001011000110: data = 6'b010101;
12'b0001011000111: data = 6'b010101;
12'b0001011001000: data = 6'b010101;
12'b0001011001001: data = 6'b010101;
12'b0001011001010: data = 6'b010101;
12'b0001011001011: data = 6'b010101;
12'b0001011001100: data = 6'b010101;
12'b0001011001101: data = 6'b010101;
12'b0001011001110: data = 6'b010101;
12'b0001011001111: data = 6'b010101;
12'b0001011010000: data = 6'b010101;
12'b0001011010001: data = 6'b010101;
12'b0001011010010: data = 6'b010101;
12'b0001011010011: data = 6'b010101;
12'b0001011010100: data = 6'b010101;
12'b0001011010101: data = 6'b010101;
12'b0001011010110: data = 6'b010101;
12'b0001011010111: data = 6'b010101;
12'b0001011011000: data = 6'b010101;
12'b0001011011001: data = 6'b010101;
12'b0001011011010: data = 6'b010101;
12'b0001011011011: data = 6'b010101;
12'b0001011011100: data = 6'b010101;
12'b0001011011101: data = 6'b010101;
12'b0001011011110: data = 6'b010101;
12'b0001011011111: data = 6'b010101;
12'b0001011100000: data = 6'b010101;
12'b0001011100001: data = 6'b010101;
12'b0001011100010: data = 6'b010101;
12'b0001011100011: data = 6'b010101;
12'b0001011100100: data = 6'b010101;
12'b0001011100101: data = 6'b010101;
12'b0001011100110: data = 6'b010101;
12'b0001011100111: data = 6'b010101;
12'b0001011101000: data = 6'b010101;
12'b0001011101001: data = 6'b010101;
12'b0001011101010: data = 6'b010101;
12'b0001011101011: data = 6'b010101;
12'b0001011101100: data = 6'b010101;
12'b0001011101101: data = 6'b010101;
12'b0001011101110: data = 6'b010101;
12'b0001011101111: data = 6'b010101;
12'b0001011110000: data = 6'b010101;
12'b0001011110001: data = 6'b010101;
12'b0001011110010: data = 6'b010101;
12'b0001011110011: data = 6'b010101;
12'b0001011110100: data = 6'b010101;
12'b0001011110101: data = 6'b010101;
12'b0001011110110: data = 6'b010101;
12'b0001011110111: data = 6'b010101;
12'b0001011111000: data = 6'b010101;
12'b0001011111001: data = 6'b010101;
12'b0001011111010: data = 6'b010101;
12'b0001011111011: data = 6'b010101;
12'b0001011111100: data = 6'b010101;
12'b0001011111101: data = 6'b010101;
12'b0001011111110: data = 6'b010101;
12'b0001011111111: data = 6'b010101;
12'b00010110000000: data = 6'b010101;
12'b00010110000001: data = 6'b010101;
12'b00010110000010: data = 6'b010101;
12'b00010110000011: data = 6'b010101;
12'b00010110000100: data = 6'b010101;
12'b00010110000101: data = 6'b010101;
12'b00010110000110: data = 6'b101010;
12'b00010110000111: data = 6'b101010;
12'b00010110001000: data = 6'b101010;
12'b00010110001001: data = 6'b101010;
12'b00010110001010: data = 6'b101010;
12'b00010110001011: data = 6'b101010;
12'b00010110001100: data = 6'b101010;
12'b00010110001101: data = 6'b101010;
12'b00010110001110: data = 6'b101010;
12'b00010110001111: data = 6'b101010;
12'b00010110010000: data = 6'b101010;
12'b00010110010001: data = 6'b010101;
12'b00010110010010: data = 6'b010101;
12'b00010110010011: data = 6'b010101;
12'b00010110010100: data = 6'b010101;
12'b00010110010101: data = 6'b010101;
12'b00010110010110: data = 6'b010101;
12'b00010110010111: data = 6'b010101;
12'b00010110011000: data = 6'b010101;
12'b00010110011001: data = 6'b010101;
12'b00010110011010: data = 6'b010101;
12'b00010110011011: data = 6'b010101;
12'b00010110011100: data = 6'b010101;
12'b00010110011101: data = 6'b010101;
12'b00010110011110: data = 6'b010101;
12'b00010110011111: data = 6'b010101;
12'b00010110100000: data = 6'b010101;
12'b00010110100001: data = 6'b010101;
12'b00010110100010: data = 6'b010101;
12'b00010110100011: data = 6'b010101;
12'b00010110100100: data = 6'b010101;
12'b00010110100101: data = 6'b010101;
12'b00010110100110: data = 6'b010101;
12'b00010110100111: data = 6'b010101;
12'b00010110101000: data = 6'b010101;
12'b00010110101001: data = 6'b010101;
12'b00010110101010: data = 6'b010101;
12'b000110000000: data = 6'b010101;
12'b000110000001: data = 6'b010101;
12'b000110000010: data = 6'b010101;
12'b000110000011: data = 6'b010101;
12'b000110000100: data = 6'b010101;
12'b000110000101: data = 6'b010101;
12'b000110000110: data = 6'b010101;
12'b000110000111: data = 6'b010101;
12'b000110001000: data = 6'b010101;
12'b000110001001: data = 6'b010101;
12'b000110001010: data = 6'b010101;
12'b000110001011: data = 6'b010101;
12'b000110001100: data = 6'b010101;
12'b000110001101: data = 6'b010101;
12'b000110001110: data = 6'b010101;
12'b000110001111: data = 6'b010101;
12'b000110010000: data = 6'b010101;
12'b000110010001: data = 6'b010101;
12'b000110010010: data = 6'b010101;
12'b000110010011: data = 6'b010101;
12'b000110010100: data = 6'b010101;
12'b000110010101: data = 6'b010101;
12'b000110010110: data = 6'b010101;
12'b000110010111: data = 6'b010101;
12'b000110011000: data = 6'b010101;
12'b000110011001: data = 6'b101010;
12'b000110011010: data = 6'b101010;
12'b000110011011: data = 6'b101010;
12'b000110011100: data = 6'b101010;
12'b000110011101: data = 6'b101010;
12'b000110011110: data = 6'b101010;
12'b000110011111: data = 6'b101010;
12'b000110100000: data = 6'b101010;
12'b000110100001: data = 6'b101010;
12'b000110100010: data = 6'b101010;
12'b000110100011: data = 6'b101010;
12'b000110100100: data = 6'b101010;
12'b000110100101: data = 6'b010101;
12'b000110100110: data = 6'b010101;
12'b000110100111: data = 6'b010101;
12'b000110101000: data = 6'b010101;
12'b000110101001: data = 6'b010101;
12'b000110101010: data = 6'b010101;
12'b000110101011: data = 6'b010101;
12'b000110101100: data = 6'b010101;
12'b000110101101: data = 6'b010101;
12'b000110101110: data = 6'b010101;
12'b000110101111: data = 6'b010101;
12'b000110110000: data = 6'b010101;
12'b000110110001: data = 6'b010101;
12'b000110110010: data = 6'b010101;
12'b000110110011: data = 6'b010101;
12'b000110110100: data = 6'b010101;
12'b000110110101: data = 6'b010101;
12'b000110110110: data = 6'b010101;
12'b000110110111: data = 6'b010101;
12'b000110111000: data = 6'b010101;
12'b000110111001: data = 6'b010101;
12'b000110111010: data = 6'b010101;
12'b000110111011: data = 6'b010101;
12'b000110111100: data = 6'b010101;
12'b000110111101: data = 6'b010101;
12'b000110111110: data = 6'b010101;
12'b000110111111: data = 6'b010101;
12'b0001101000000: data = 6'b010101;
12'b0001101000001: data = 6'b010101;
12'b0001101000010: data = 6'b010101;
12'b0001101000011: data = 6'b010101;
12'b0001101000100: data = 6'b010101;
12'b0001101000101: data = 6'b010101;
12'b0001101000110: data = 6'b010101;
12'b0001101000111: data = 6'b010101;
12'b0001101001000: data = 6'b010101;
12'b0001101001001: data = 6'b010101;
12'b0001101001010: data = 6'b010101;
12'b0001101001011: data = 6'b010101;
12'b0001101001100: data = 6'b010101;
12'b0001101001101: data = 6'b010101;
12'b0001101001110: data = 6'b010101;
12'b0001101001111: data = 6'b010101;
12'b0001101010000: data = 6'b010101;
12'b0001101010001: data = 6'b010101;
12'b0001101010010: data = 6'b010101;
12'b0001101010011: data = 6'b010101;
12'b0001101010100: data = 6'b010101;
12'b0001101010101: data = 6'b010101;
12'b0001101010110: data = 6'b010101;
12'b0001101010111: data = 6'b010101;
12'b0001101011000: data = 6'b010101;
12'b0001101011001: data = 6'b010101;
12'b0001101011010: data = 6'b010101;
12'b0001101011011: data = 6'b010101;
12'b0001101011100: data = 6'b010101;
12'b0001101011101: data = 6'b010101;
12'b0001101011110: data = 6'b010101;
12'b0001101011111: data = 6'b010101;
12'b0001101100000: data = 6'b010101;
12'b0001101100001: data = 6'b010101;
12'b0001101100010: data = 6'b010101;
12'b0001101100011: data = 6'b010101;
12'b0001101100100: data = 6'b010101;
12'b0001101100101: data = 6'b010101;
12'b0001101100110: data = 6'b010101;
12'b0001101100111: data = 6'b010101;
12'b0001101101000: data = 6'b010101;
12'b0001101101001: data = 6'b010101;
12'b0001101101010: data = 6'b010101;
12'b0001101101011: data = 6'b010101;
12'b0001101101100: data = 6'b010101;
12'b0001101101101: data = 6'b010101;
12'b0001101101110: data = 6'b010101;
12'b0001101101111: data = 6'b010101;
12'b0001101110000: data = 6'b010101;
12'b0001101110001: data = 6'b010101;
12'b0001101110010: data = 6'b010101;
12'b0001101110011: data = 6'b010101;
12'b0001101110100: data = 6'b010101;
12'b0001101110101: data = 6'b010101;
12'b0001101110110: data = 6'b010101;
12'b0001101110111: data = 6'b010101;
12'b0001101111000: data = 6'b010101;
12'b0001101111001: data = 6'b010101;
12'b0001101111010: data = 6'b010101;
12'b0001101111011: data = 6'b010101;
12'b0001101111100: data = 6'b010101;
12'b0001101111101: data = 6'b010101;
12'b0001101111110: data = 6'b010101;
12'b0001101111111: data = 6'b010101;
12'b00011010000000: data = 6'b010101;
12'b00011010000001: data = 6'b010101;
12'b00011010000010: data = 6'b010101;
12'b00011010000011: data = 6'b010101;
12'b00011010000100: data = 6'b010101;
12'b00011010000101: data = 6'b010101;
12'b00011010000110: data = 6'b101010;
12'b00011010000111: data = 6'b101010;
12'b00011010001000: data = 6'b101010;
12'b00011010001001: data = 6'b101010;
12'b00011010001010: data = 6'b101010;
12'b00011010001011: data = 6'b101010;
12'b00011010001100: data = 6'b111111;
12'b00011010001101: data = 6'b101010;
12'b00011010001110: data = 6'b101010;
12'b00011010001111: data = 6'b101010;
12'b00011010010000: data = 6'b101010;
12'b00011010010001: data = 6'b101010;
12'b00011010010010: data = 6'b010101;
12'b00011010010011: data = 6'b010101;
12'b00011010010100: data = 6'b010101;
12'b00011010010101: data = 6'b010101;
12'b00011010010110: data = 6'b010101;
12'b00011010010111: data = 6'b010101;
12'b00011010011000: data = 6'b010101;
12'b00011010011001: data = 6'b010101;
12'b00011010011010: data = 6'b010101;
12'b00011010011011: data = 6'b010101;
12'b00011010011100: data = 6'b010101;
12'b00011010011101: data = 6'b010101;
12'b00011010011110: data = 6'b010101;
12'b00011010011111: data = 6'b010101;
12'b00011010100000: data = 6'b010101;
12'b00011010100001: data = 6'b010101;
12'b00011010100010: data = 6'b010101;
12'b00011010100011: data = 6'b010101;
12'b00011010100100: data = 6'b010101;
12'b00011010100101: data = 6'b010101;
12'b00011010100110: data = 6'b010101;
12'b00011010100111: data = 6'b010101;
12'b00011010101000: data = 6'b010101;
12'b00011010101001: data = 6'b010101;
12'b00011010101010: data = 6'b010101;
12'b000111000000: data = 6'b010101;
12'b000111000001: data = 6'b010101;
12'b000111000010: data = 6'b010101;
12'b000111000011: data = 6'b010101;
12'b000111000100: data = 6'b010101;
12'b000111000101: data = 6'b010101;
12'b000111000110: data = 6'b010101;
12'b000111000111: data = 6'b010101;
12'b000111001000: data = 6'b010101;
12'b000111001001: data = 6'b010101;
12'b000111001010: data = 6'b010101;
12'b000111001011: data = 6'b010101;
12'b000111001100: data = 6'b010101;
12'b000111001101: data = 6'b010101;
12'b000111001110: data = 6'b010101;
12'b000111001111: data = 6'b010101;
12'b000111010000: data = 6'b010101;
12'b000111010001: data = 6'b010101;
12'b000111010010: data = 6'b010101;
12'b000111010011: data = 6'b010101;
12'b000111010100: data = 6'b010101;
12'b000111010101: data = 6'b010101;
12'b000111010110: data = 6'b010101;
12'b000111010111: data = 6'b010101;
12'b000111011000: data = 6'b010101;
12'b000111011001: data = 6'b101010;
12'b000111011010: data = 6'b101010;
12'b000111011011: data = 6'b101010;
12'b000111011100: data = 6'b101010;
12'b000111011101: data = 6'b101010;
12'b000111011110: data = 6'b101010;
12'b000111011111: data = 6'b101010;
12'b000111100000: data = 6'b101010;
12'b000111100001: data = 6'b101010;
12'b000111100010: data = 6'b101010;
12'b000111100011: data = 6'b101010;
12'b000111100100: data = 6'b101010;
12'b000111100101: data = 6'b010101;
12'b000111100110: data = 6'b010101;
12'b000111100111: data = 6'b010101;
12'b000111101000: data = 6'b010101;
12'b000111101001: data = 6'b010101;
12'b000111101010: data = 6'b010101;
12'b000111101011: data = 6'b010101;
12'b000111101100: data = 6'b010101;
12'b000111101101: data = 6'b010101;
12'b000111101110: data = 6'b010101;
12'b000111101111: data = 6'b010101;
12'b000111110000: data = 6'b010101;
12'b000111110001: data = 6'b010101;
12'b000111110010: data = 6'b010101;
12'b000111110011: data = 6'b010101;
12'b000111110100: data = 6'b010101;
12'b000111110101: data = 6'b010101;
12'b000111110110: data = 6'b010101;
12'b000111110111: data = 6'b010101;
12'b000111111000: data = 6'b010101;
12'b000111111001: data = 6'b100101;
12'b000111111010: data = 6'b100101;
12'b000111111011: data = 6'b100101;
12'b000111111100: data = 6'b100101;
12'b000111111101: data = 6'b100101;
12'b000111111110: data = 6'b100101;
12'b000111111111: data = 6'b100101;
12'b0001111000000: data = 6'b100101;
12'b0001111000001: data = 6'b100101;
12'b0001111000010: data = 6'b100101;
12'b0001111000011: data = 6'b100101;
12'b0001111000100: data = 6'b100101;
12'b0001111000101: data = 6'b100101;
12'b0001111000110: data = 6'b100101;
12'b0001111000111: data = 6'b100101;
12'b0001111001000: data = 6'b100101;
12'b0001111001001: data = 6'b100101;
12'b0001111001010: data = 6'b100101;
12'b0001111001011: data = 6'b100101;
12'b0001111001100: data = 6'b100101;
12'b0001111001101: data = 6'b100101;
12'b0001111001110: data = 6'b100101;
12'b0001111001111: data = 6'b100101;
12'b0001111010000: data = 6'b100101;
12'b0001111010001: data = 6'b100101;
12'b0001111010010: data = 6'b100101;
12'b0001111010011: data = 6'b100101;
12'b0001111010100: data = 6'b100101;
12'b0001111010101: data = 6'b010101;
12'b0001111010110: data = 6'b010101;
12'b0001111010111: data = 6'b010101;
12'b0001111011000: data = 6'b010101;
12'b0001111011001: data = 6'b010101;
12'b0001111011010: data = 6'b010101;
12'b0001111011011: data = 6'b010101;
12'b0001111011100: data = 6'b010101;
12'b0001111011101: data = 6'b010101;
12'b0001111011110: data = 6'b010101;
12'b0001111011111: data = 6'b010101;
12'b0001111100000: data = 6'b010101;
12'b0001111100001: data = 6'b010101;
12'b0001111100010: data = 6'b010101;
12'b0001111100011: data = 6'b010101;
12'b0001111100100: data = 6'b010101;
12'b0001111100101: data = 6'b010101;
12'b0001111100110: data = 6'b010101;
12'b0001111100111: data = 6'b010101;
12'b0001111101000: data = 6'b010101;
12'b0001111101001: data = 6'b010101;
12'b0001111101010: data = 6'b010101;
12'b0001111101011: data = 6'b010101;
12'b0001111101100: data = 6'b010101;
12'b0001111101101: data = 6'b010101;
12'b0001111101110: data = 6'b010101;
12'b0001111101111: data = 6'b010101;
12'b0001111110000: data = 6'b010101;
12'b0001111110001: data = 6'b010101;
12'b0001111110010: data = 6'b010101;
12'b0001111110011: data = 6'b010101;
12'b0001111110100: data = 6'b010101;
12'b0001111110101: data = 6'b010101;
12'b0001111110110: data = 6'b010101;
12'b0001111110111: data = 6'b010101;
12'b0001111111000: data = 6'b010101;
12'b0001111111001: data = 6'b010101;
12'b0001111111010: data = 6'b010101;
12'b0001111111011: data = 6'b010101;
12'b0001111111100: data = 6'b010101;
12'b0001111111101: data = 6'b010101;
12'b0001111111110: data = 6'b010101;
12'b0001111111111: data = 6'b010101;
12'b00011110000000: data = 6'b010101;
12'b00011110000001: data = 6'b010101;
12'b00011110000010: data = 6'b010101;
12'b00011110000011: data = 6'b010101;
12'b00011110000100: data = 6'b010101;
12'b00011110000101: data = 6'b010101;
12'b00011110000110: data = 6'b101001;
12'b00011110000111: data = 6'b101010;
12'b00011110001000: data = 6'b101010;
12'b00011110001001: data = 6'b101010;
12'b00011110001010: data = 6'b101010;
12'b00011110001011: data = 6'b101010;
12'b00011110001100: data = 6'b101010;
12'b00011110001101: data = 6'b101010;
12'b00011110001110: data = 6'b101010;
12'b00011110001111: data = 6'b101010;
12'b00011110010000: data = 6'b101010;
12'b00011110010001: data = 6'b101010;
12'b00011110010010: data = 6'b010101;
12'b00011110010011: data = 6'b010101;
12'b00011110010100: data = 6'b010101;
12'b00011110010101: data = 6'b010101;
12'b00011110010110: data = 6'b010101;
12'b00011110010111: data = 6'b010101;
12'b00011110011000: data = 6'b010101;
12'b00011110011001: data = 6'b010101;
12'b00011110011010: data = 6'b010101;
12'b00011110011011: data = 6'b010101;
12'b00011110011100: data = 6'b010101;
12'b00011110011101: data = 6'b010101;
12'b00011110011110: data = 6'b010101;
12'b00011110011111: data = 6'b010101;
12'b00011110100000: data = 6'b010101;
12'b00011110100001: data = 6'b010101;
12'b00011110100010: data = 6'b010101;
12'b00011110100011: data = 6'b010101;
12'b00011110100100: data = 6'b010101;
12'b00011110100101: data = 6'b010101;
12'b00011110100110: data = 6'b010101;
12'b00011110100111: data = 6'b010101;
12'b00011110101000: data = 6'b010101;
12'b00011110101001: data = 6'b010101;
12'b00011110101010: data = 6'b010101;
12'b001000000000: data = 6'b010101;
12'b001000000001: data = 6'b010101;
12'b001000000010: data = 6'b010101;
12'b001000000011: data = 6'b010101;
12'b001000000100: data = 6'b010101;
12'b001000000101: data = 6'b010101;
12'b001000000110: data = 6'b010101;
12'b001000000111: data = 6'b010101;
12'b001000001000: data = 6'b010101;
12'b001000001001: data = 6'b010101;
12'b001000001010: data = 6'b010101;
12'b001000001011: data = 6'b010101;
12'b001000001100: data = 6'b010101;
12'b001000001101: data = 6'b010101;
12'b001000001110: data = 6'b010101;
12'b001000001111: data = 6'b010101;
12'b001000010000: data = 6'b010101;
12'b001000010001: data = 6'b010101;
12'b001000010010: data = 6'b010101;
12'b001000010011: data = 6'b010101;
12'b001000010100: data = 6'b010101;
12'b001000010101: data = 6'b010101;
12'b001000010110: data = 6'b010101;
12'b001000010111: data = 6'b010101;
12'b001000011000: data = 6'b010101;
12'b001000011001: data = 6'b101010;
12'b001000011010: data = 6'b101010;
12'b001000011011: data = 6'b101010;
12'b001000011100: data = 6'b010101;
12'b001000011101: data = 6'b000000;
12'b001000011110: data = 6'b000000;
12'b001000011111: data = 6'b010101;
12'b001000100000: data = 6'b010101;
12'b001000100001: data = 6'b010101;
12'b001000100010: data = 6'b010101;
12'b001000100011: data = 6'b010101;
12'b001000100100: data = 6'b010101;
12'b001000100101: data = 6'b010101;
12'b001000100110: data = 6'b010101;
12'b001000100111: data = 6'b010101;
12'b001000101000: data = 6'b101001;
12'b001000101001: data = 6'b101001;
12'b001000101010: data = 6'b101010;
12'b001000101011: data = 6'b101010;
12'b001000101100: data = 6'b101010;
12'b001000101101: data = 6'b101010;
12'b001000101110: data = 6'b101010;
12'b001000101111: data = 6'b101010;
12'b001000110000: data = 6'b101010;
12'b001000110001: data = 6'b101010;
12'b001000110010: data = 6'b101010;
12'b001000110011: data = 6'b101010;
12'b001000110100: data = 6'b101010;
12'b001000110101: data = 6'b101010;
12'b001000110110: data = 6'b101010;
12'b001000110111: data = 6'b101010;
12'b001000111000: data = 6'b101010;
12'b001000111001: data = 6'b111111;
12'b001000111010: data = 6'b111111;
12'b001000111011: data = 6'b111111;
12'b001000111100: data = 6'b111111;
12'b001000111101: data = 6'b111111;
12'b001000111110: data = 6'b111111;
12'b001000111111: data = 6'b111111;
12'b0010001000000: data = 6'b111111;
12'b0010001000001: data = 6'b111111;
12'b0010001000010: data = 6'b111111;
12'b0010001000011: data = 6'b111111;
12'b0010001000100: data = 6'b111111;
12'b0010001000101: data = 6'b111111;
12'b0010001000110: data = 6'b111111;
12'b0010001000111: data = 6'b111111;
12'b0010001001000: data = 6'b111111;
12'b0010001001001: data = 6'b111111;
12'b0010001001010: data = 6'b111111;
12'b0010001001011: data = 6'b111111;
12'b0010001001100: data = 6'b111111;
12'b0010001001101: data = 6'b111110;
12'b0010001001110: data = 6'b111110;
12'b0010001001111: data = 6'b111110;
12'b0010001010000: data = 6'b111110;
12'b0010001010001: data = 6'b101010;
12'b0010001010010: data = 6'b101010;
12'b0010001010011: data = 6'b101010;
12'b0010001010100: data = 6'b101010;
12'b0010001010101: data = 6'b101010;
12'b0010001010110: data = 6'b101010;
12'b0010001010111: data = 6'b101010;
12'b0010001011000: data = 6'b101010;
12'b0010001011001: data = 6'b101010;
12'b0010001011010: data = 6'b101010;
12'b0010001011011: data = 6'b101010;
12'b0010001011100: data = 6'b101010;
12'b0010001011101: data = 6'b101010;
12'b0010001011110: data = 6'b101010;
12'b0010001011111: data = 6'b101010;
12'b0010001100000: data = 6'b101010;
12'b0010001100001: data = 6'b101010;
12'b0010001100010: data = 6'b101010;
12'b0010001100011: data = 6'b101010;
12'b0010001100100: data = 6'b101010;
12'b0010001100101: data = 6'b101010;
12'b0010001100110: data = 6'b101010;
12'b0010001100111: data = 6'b101010;
12'b0010001101000: data = 6'b101010;
12'b0010001101001: data = 6'b101010;
12'b0010001101010: data = 6'b101010;
12'b0010001101011: data = 6'b101010;
12'b0010001101100: data = 6'b101010;
12'b0010001101101: data = 6'b101010;
12'b0010001101110: data = 6'b101010;
12'b0010001101111: data = 6'b101010;
12'b0010001110000: data = 6'b101010;
12'b0010001110001: data = 6'b101010;
12'b0010001110010: data = 6'b101010;
12'b0010001110011: data = 6'b101010;
12'b0010001110100: data = 6'b101001;
12'b0010001110101: data = 6'b101001;
12'b0010001110110: data = 6'b010101;
12'b0010001110111: data = 6'b010101;
12'b0010001111000: data = 6'b010101;
12'b0010001111001: data = 6'b010101;
12'b0010001111010: data = 6'b010101;
12'b0010001111011: data = 6'b010101;
12'b0010001111100: data = 6'b010101;
12'b0010001111101: data = 6'b010101;
12'b0010001111110: data = 6'b010101;
12'b0010001111111: data = 6'b010101;
12'b00100010000000: data = 6'b010101;
12'b00100010000001: data = 6'b010101;
12'b00100010000010: data = 6'b010101;
12'b00100010000011: data = 6'b010101;
12'b00100010000100: data = 6'b010101;
12'b00100010000101: data = 6'b010101;
12'b00100010000110: data = 6'b010101;
12'b00100010000111: data = 6'b010101;
12'b00100010001000: data = 6'b010101;
12'b00100010001001: data = 6'b010101;
12'b00100010001010: data = 6'b010101;
12'b00100010001011: data = 6'b010101;
12'b00100010001100: data = 6'b000000;
12'b00100010001101: data = 6'b010101;
12'b00100010001110: data = 6'b101010;
12'b00100010001111: data = 6'b101010;
12'b00100010010000: data = 6'b101010;
12'b00100010010001: data = 6'b101010;
12'b00100010010010: data = 6'b010101;
12'b00100010010011: data = 6'b010101;
12'b00100010010100: data = 6'b010101;
12'b00100010010101: data = 6'b010101;
12'b00100010010110: data = 6'b010101;
12'b00100010010111: data = 6'b010101;
12'b00100010011000: data = 6'b010101;
12'b00100010011001: data = 6'b010101;
12'b00100010011010: data = 6'b010101;
12'b00100010011011: data = 6'b010101;
12'b00100010011100: data = 6'b010101;
12'b00100010011101: data = 6'b010101;
12'b00100010011110: data = 6'b010101;
12'b00100010011111: data = 6'b010101;
12'b00100010100000: data = 6'b010101;
12'b00100010100001: data = 6'b010101;
12'b00100010100010: data = 6'b010101;
12'b00100010100011: data = 6'b010101;
12'b00100010100100: data = 6'b010101;
12'b00100010100101: data = 6'b010101;
12'b00100010100110: data = 6'b010101;
12'b00100010100111: data = 6'b010101;
12'b00100010101000: data = 6'b010101;
12'b00100010101001: data = 6'b010101;
12'b00100010101010: data = 6'b010101;
12'b001001000000: data = 6'b010101;
12'b001001000001: data = 6'b010101;
12'b001001000010: data = 6'b010101;
12'b001001000011: data = 6'b010101;
12'b001001000100: data = 6'b010101;
12'b001001000101: data = 6'b010101;
12'b001001000110: data = 6'b010101;
12'b001001000111: data = 6'b010101;
12'b001001001000: data = 6'b010101;
12'b001001001001: data = 6'b010101;
12'b001001001010: data = 6'b010101;
12'b001001001011: data = 6'b010101;
12'b001001001100: data = 6'b010101;
12'b001001001101: data = 6'b010101;
12'b001001001110: data = 6'b010101;
12'b001001001111: data = 6'b010101;
12'b001001010000: data = 6'b010101;
12'b001001010001: data = 6'b010101;
12'b001001010010: data = 6'b010101;
12'b001001010011: data = 6'b010101;
12'b001001010100: data = 6'b010101;
12'b001001010101: data = 6'b010101;
12'b001001010110: data = 6'b010101;
12'b001001010111: data = 6'b010101;
12'b001001011000: data = 6'b010101;
12'b001001011001: data = 6'b101010;
12'b001001011010: data = 6'b101010;
12'b001001011011: data = 6'b101010;
12'b001001011100: data = 6'b010101;
12'b001001011101: data = 6'b000000;
12'b001001011110: data = 6'b000000;
12'b001001011111: data = 6'b000000;
12'b001001100000: data = 6'b010101;
12'b001001100001: data = 6'b010101;
12'b001001100010: data = 6'b010101;
12'b001001100011: data = 6'b010101;
12'b001001100100: data = 6'b010101;
12'b001001100101: data = 6'b010101;
12'b001001100110: data = 6'b010101;
12'b001001100111: data = 6'b010101;
12'b001001101000: data = 6'b101001;
12'b001001101001: data = 6'b101001;
12'b001001101010: data = 6'b101010;
12'b001001101011: data = 6'b101010;
12'b001001101100: data = 6'b101010;
12'b001001101101: data = 6'b101010;
12'b001001101110: data = 6'b101010;
12'b001001101111: data = 6'b101010;
12'b001001110000: data = 6'b101010;
12'b001001110001: data = 6'b101010;
12'b001001110010: data = 6'b101010;
12'b001001110011: data = 6'b101010;
12'b001001110100: data = 6'b101010;
12'b001001110101: data = 6'b101010;
12'b001001110110: data = 6'b101010;
12'b001001110111: data = 6'b111111;
12'b001001111000: data = 6'b111111;
12'b001001111001: data = 6'b111111;
12'b001001111010: data = 6'b111111;
12'b001001111011: data = 6'b111111;
12'b001001111100: data = 6'b111111;
12'b001001111101: data = 6'b111111;
12'b001001111110: data = 6'b111111;
12'b001001111111: data = 6'b111111;
12'b0010011000000: data = 6'b111111;
12'b0010011000001: data = 6'b111111;
12'b0010011000010: data = 6'b111111;
12'b0010011000011: data = 6'b111111;
12'b0010011000100: data = 6'b111111;
12'b0010011000101: data = 6'b111111;
12'b0010011000110: data = 6'b111111;
12'b0010011000111: data = 6'b111111;
12'b0010011001000: data = 6'b111111;
12'b0010011001001: data = 6'b111111;
12'b0010011001010: data = 6'b111111;
12'b0010011001011: data = 6'b111111;
12'b0010011001100: data = 6'b111111;
12'b0010011001101: data = 6'b111111;
12'b0010011001110: data = 6'b111111;
12'b0010011001111: data = 6'b111111;
12'b0010011010000: data = 6'b111111;
12'b0010011010001: data = 6'b111110;
12'b0010011010010: data = 6'b111111;
12'b0010011010011: data = 6'b111110;
12'b0010011010100: data = 6'b111111;
12'b0010011010101: data = 6'b111110;
12'b0010011010110: data = 6'b111110;
12'b0010011010111: data = 6'b101010;
12'b0010011011000: data = 6'b101010;
12'b0010011011001: data = 6'b101010;
12'b0010011011010: data = 6'b101010;
12'b0010011011011: data = 6'b101010;
12'b0010011011100: data = 6'b101010;
12'b0010011011101: data = 6'b101010;
12'b0010011011110: data = 6'b101010;
12'b0010011011111: data = 6'b101010;
12'b0010011100000: data = 6'b101010;
12'b0010011100001: data = 6'b101010;
12'b0010011100010: data = 6'b101010;
12'b0010011100011: data = 6'b101010;
12'b0010011100100: data = 6'b101010;
12'b0010011100101: data = 6'b101010;
12'b0010011100110: data = 6'b101010;
12'b0010011100111: data = 6'b101010;
12'b0010011101000: data = 6'b101010;
12'b0010011101001: data = 6'b101010;
12'b0010011101010: data = 6'b101010;
12'b0010011101011: data = 6'b101010;
12'b0010011101100: data = 6'b101010;
12'b0010011101101: data = 6'b101010;
12'b0010011101110: data = 6'b101010;
12'b0010011101111: data = 6'b101010;
12'b0010011110000: data = 6'b101010;
12'b0010011110001: data = 6'b101010;
12'b0010011110010: data = 6'b101010;
12'b0010011110011: data = 6'b101010;
12'b0010011110100: data = 6'b101001;
12'b0010011110101: data = 6'b101001;
12'b0010011110110: data = 6'b010101;
12'b0010011110111: data = 6'b010101;
12'b0010011111000: data = 6'b010101;
12'b0010011111001: data = 6'b010101;
12'b0010011111010: data = 6'b010101;
12'b0010011111011: data = 6'b010101;
12'b0010011111100: data = 6'b010101;
12'b0010011111101: data = 6'b010101;
12'b0010011111110: data = 6'b010101;
12'b0010011111111: data = 6'b010101;
12'b00100110000000: data = 6'b010101;
12'b00100110000001: data = 6'b010101;
12'b00100110000010: data = 6'b010101;
12'b00100110000011: data = 6'b010101;
12'b00100110000100: data = 6'b010101;
12'b00100110000101: data = 6'b010101;
12'b00100110000110: data = 6'b010101;
12'b00100110000111: data = 6'b010101;
12'b00100110001000: data = 6'b010101;
12'b00100110001001: data = 6'b010101;
12'b00100110001010: data = 6'b010101;
12'b00100110001011: data = 6'b010101;
12'b00100110001100: data = 6'b000000;
12'b00100110001101: data = 6'b000000;
12'b00100110001110: data = 6'b101010;
12'b00100110001111: data = 6'b101010;
12'b00100110010000: data = 6'b101010;
12'b00100110010001: data = 6'b101010;
12'b00100110010010: data = 6'b010101;
12'b00100110010011: data = 6'b010101;
12'b00100110010100: data = 6'b010101;
12'b00100110010101: data = 6'b010101;
12'b00100110010110: data = 6'b010101;
12'b00100110010111: data = 6'b010101;
12'b00100110011000: data = 6'b010101;
12'b00100110011001: data = 6'b010101;
12'b00100110011010: data = 6'b010101;
12'b00100110011011: data = 6'b010101;
12'b00100110011100: data = 6'b010101;
12'b00100110011101: data = 6'b010101;
12'b00100110011110: data = 6'b010101;
12'b00100110011111: data = 6'b010101;
12'b00100110100000: data = 6'b010101;
12'b00100110100001: data = 6'b010101;
12'b00100110100010: data = 6'b010101;
12'b00100110100011: data = 6'b010101;
12'b00100110100100: data = 6'b010101;
12'b00100110100101: data = 6'b010101;
12'b00100110100110: data = 6'b010101;
12'b00100110100111: data = 6'b010101;
12'b00100110101000: data = 6'b010101;
12'b00100110101001: data = 6'b010101;
12'b00100110101010: data = 6'b010101;
12'b001010000000: data = 6'b010101;
12'b001010000001: data = 6'b010101;
12'b001010000010: data = 6'b010101;
12'b001010000011: data = 6'b010101;
12'b001010000100: data = 6'b010101;
12'b001010000101: data = 6'b010101;
12'b001010000110: data = 6'b010101;
12'b001010000111: data = 6'b010101;
12'b001010001000: data = 6'b010101;
12'b001010001001: data = 6'b010101;
12'b001010001010: data = 6'b010101;
12'b001010001011: data = 6'b010101;
12'b001010001100: data = 6'b010101;
12'b001010001101: data = 6'b010101;
12'b001010001110: data = 6'b010101;
12'b001010001111: data = 6'b010101;
12'b001010010000: data = 6'b010101;
12'b001010010001: data = 6'b010101;
12'b001010010010: data = 6'b010101;
12'b001010010011: data = 6'b010101;
12'b001010010100: data = 6'b010101;
12'b001010010101: data = 6'b010101;
12'b001010010110: data = 6'b010101;
12'b001010010111: data = 6'b010101;
12'b001010011000: data = 6'b010101;
12'b001010011001: data = 6'b101010;
12'b001010011010: data = 6'b101010;
12'b001010011011: data = 6'b101010;
12'b001010011100: data = 6'b010101;
12'b001010011101: data = 6'b000000;
12'b001010011110: data = 6'b000000;
12'b001010011111: data = 6'b010101;
12'b001010100000: data = 6'b101010;
12'b001010100001: data = 6'b101010;
12'b001010100010: data = 6'b101010;
12'b001010100011: data = 6'b101010;
12'b001010100100: data = 6'b101010;
12'b001010100101: data = 6'b101010;
12'b001010100110: data = 6'b101010;
12'b001010100111: data = 6'b101010;
12'b001010101000: data = 6'b101010;
12'b001010101001: data = 6'b101010;
12'b001010101010: data = 6'b101010;
12'b001010101011: data = 6'b101010;
12'b001010101100: data = 6'b101010;
12'b001010101101: data = 6'b101010;
12'b001010101110: data = 6'b101010;
12'b001010101111: data = 6'b101010;
12'b001010110000: data = 6'b101010;
12'b001010110001: data = 6'b101010;
12'b001010110010: data = 6'b101010;
12'b001010110011: data = 6'b101010;
12'b001010110100: data = 6'b111010;
12'b001010110101: data = 6'b111110;
12'b001010110110: data = 6'b111110;
12'b001010110111: data = 6'b111111;
12'b001010111000: data = 6'b111111;
12'b001010111001: data = 6'b111111;
12'b001010111010: data = 6'b111111;
12'b001010111011: data = 6'b111111;
12'b001010111100: data = 6'b111111;
12'b001010111101: data = 6'b111111;
12'b001010111110: data = 6'b111111;
12'b001010111111: data = 6'b111111;
12'b0010101000000: data = 6'b111111;
12'b0010101000001: data = 6'b111111;
12'b0010101000010: data = 6'b111111;
12'b0010101000011: data = 6'b111111;
12'b0010101000100: data = 6'b111111;
12'b0010101000101: data = 6'b111111;
12'b0010101000110: data = 6'b111111;
12'b0010101000111: data = 6'b111111;
12'b0010101001000: data = 6'b111111;
12'b0010101001001: data = 6'b111111;
12'b0010101001010: data = 6'b111111;
12'b0010101001011: data = 6'b111111;
12'b0010101001100: data = 6'b111111;
12'b0010101001101: data = 6'b111111;
12'b0010101001110: data = 6'b111111;
12'b0010101001111: data = 6'b111111;
12'b0010101010000: data = 6'b111111;
12'b0010101010001: data = 6'b111111;
12'b0010101010010: data = 6'b111111;
12'b0010101010011: data = 6'b111111;
12'b0010101010100: data = 6'b111110;
12'b0010101010101: data = 6'b111110;
12'b0010101010110: data = 6'b111110;
12'b0010101010111: data = 6'b111111;
12'b0010101011000: data = 6'b111111;
12'b0010101011001: data = 6'b111110;
12'b0010101011010: data = 6'b111010;
12'b0010101011011: data = 6'b111010;
12'b0010101011100: data = 6'b101010;
12'b0010101011101: data = 6'b101010;
12'b0010101011110: data = 6'b101010;
12'b0010101011111: data = 6'b101010;
12'b0010101100000: data = 6'b101010;
12'b0010101100001: data = 6'b101010;
12'b0010101100010: data = 6'b101010;
12'b0010101100011: data = 6'b101010;
12'b0010101100100: data = 6'b101010;
12'b0010101100101: data = 6'b101010;
12'b0010101100110: data = 6'b101010;
12'b0010101100111: data = 6'b101010;
12'b0010101101000: data = 6'b101010;
12'b0010101101001: data = 6'b101010;
12'b0010101101010: data = 6'b101010;
12'b0010101101011: data = 6'b101010;
12'b0010101101100: data = 6'b101010;
12'b0010101101101: data = 6'b101010;
12'b0010101101110: data = 6'b101010;
12'b0010101101111: data = 6'b101010;
12'b0010101110000: data = 6'b101010;
12'b0010101110001: data = 6'b101010;
12'b0010101110010: data = 6'b101010;
12'b0010101110011: data = 6'b101010;
12'b0010101110100: data = 6'b101010;
12'b0010101110101: data = 6'b101010;
12'b0010101110110: data = 6'b101010;
12'b0010101110111: data = 6'b101010;
12'b0010101111000: data = 6'b101010;
12'b0010101111001: data = 6'b101010;
12'b0010101111010: data = 6'b101010;
12'b0010101111011: data = 6'b101010;
12'b0010101111100: data = 6'b101010;
12'b0010101111101: data = 6'b101010;
12'b0010101111110: data = 6'b101010;
12'b0010101111111: data = 6'b101010;
12'b00101010000000: data = 6'b101010;
12'b00101010000001: data = 6'b101010;
12'b00101010000010: data = 6'b101010;
12'b00101010000011: data = 6'b101010;
12'b00101010000100: data = 6'b101010;
12'b00101010000101: data = 6'b101010;
12'b00101010000110: data = 6'b101010;
12'b00101010000111: data = 6'b101010;
12'b00101010001000: data = 6'b101010;
12'b00101010001001: data = 6'b101010;
12'b00101010001010: data = 6'b101010;
12'b00101010001011: data = 6'b010101;
12'b00101010001100: data = 6'b000000;
12'b00101010001101: data = 6'b000000;
12'b00101010001110: data = 6'b101010;
12'b00101010001111: data = 6'b101010;
12'b00101010010000: data = 6'b101010;
12'b00101010010001: data = 6'b101010;
12'b00101010010010: data = 6'b010101;
12'b00101010010011: data = 6'b010101;
12'b00101010010100: data = 6'b010101;
12'b00101010010101: data = 6'b010101;
12'b00101010010110: data = 6'b010101;
12'b00101010010111: data = 6'b010101;
12'b00101010011000: data = 6'b010101;
12'b00101010011001: data = 6'b010101;
12'b00101010011010: data = 6'b010101;
12'b00101010011011: data = 6'b010101;
12'b00101010011100: data = 6'b010101;
12'b00101010011101: data = 6'b010101;
12'b00101010011110: data = 6'b010101;
12'b00101010011111: data = 6'b010101;
12'b00101010100000: data = 6'b010101;
12'b00101010100001: data = 6'b010101;
12'b00101010100010: data = 6'b010101;
12'b00101010100011: data = 6'b010101;
12'b00101010100100: data = 6'b010101;
12'b00101010100101: data = 6'b010101;
12'b00101010100110: data = 6'b010101;
12'b00101010100111: data = 6'b010101;
12'b00101010101000: data = 6'b010101;
12'b00101010101001: data = 6'b010101;
12'b00101010101010: data = 6'b010101;
12'b001011000000: data = 6'b010101;
12'b001011000001: data = 6'b010101;
12'b001011000010: data = 6'b010101;
12'b001011000011: data = 6'b010101;
12'b001011000100: data = 6'b010101;
12'b001011000101: data = 6'b010101;
12'b001011000110: data = 6'b010101;
12'b001011000111: data = 6'b010101;
12'b001011001000: data = 6'b010101;
12'b001011001001: data = 6'b010101;
12'b001011001010: data = 6'b010101;
12'b001011001011: data = 6'b010101;
12'b001011001100: data = 6'b010101;
12'b001011001101: data = 6'b010101;
12'b001011001110: data = 6'b010101;
12'b001011001111: data = 6'b010101;
12'b001011010000: data = 6'b010101;
12'b001011010001: data = 6'b010101;
12'b001011010010: data = 6'b010101;
12'b001011010011: data = 6'b010101;
12'b001011010100: data = 6'b010101;
12'b001011010101: data = 6'b010101;
12'b001011010110: data = 6'b010101;
12'b001011010111: data = 6'b010101;
12'b001011011000: data = 6'b010101;
12'b001011011001: data = 6'b101010;
12'b001011011010: data = 6'b101010;
12'b001011011011: data = 6'b101010;
12'b001011011100: data = 6'b010101;
12'b001011011101: data = 6'b000000;
12'b001011011110: data = 6'b000000;
12'b001011011111: data = 6'b010101;
12'b001011100000: data = 6'b111111;
12'b001011100001: data = 6'b111111;
12'b001011100010: data = 6'b111111;
12'b001011100011: data = 6'b111111;
12'b001011100100: data = 6'b111111;
12'b001011100101: data = 6'b111111;
12'b001011100110: data = 6'b111111;
12'b001011100111: data = 6'b111111;
12'b001011101000: data = 6'b111111;
12'b001011101001: data = 6'b111111;
12'b001011101010: data = 6'b111111;
12'b001011101011: data = 6'b111111;
12'b001011101100: data = 6'b111111;
12'b001011101101: data = 6'b111111;
12'b001011101110: data = 6'b111111;
12'b001011101111: data = 6'b111111;
12'b001011110000: data = 6'b111111;
12'b001011110001: data = 6'b111111;
12'b001011110010: data = 6'b111111;
12'b001011110011: data = 6'b111111;
12'b001011110100: data = 6'b111111;
12'b001011110101: data = 6'b111111;
12'b001011110110: data = 6'b111111;
12'b001011110111: data = 6'b111111;
12'b001011111000: data = 6'b111111;
12'b001011111001: data = 6'b111111;
12'b001011111010: data = 6'b111111;
12'b001011111011: data = 6'b111111;
12'b001011111100: data = 6'b111111;
12'b001011111101: data = 6'b111111;
12'b001011111110: data = 6'b111111;
12'b001011111111: data = 6'b111111;
12'b0010111000000: data = 6'b111111;
12'b0010111000001: data = 6'b111111;
12'b0010111000010: data = 6'b111111;
12'b0010111000011: data = 6'b111111;
12'b0010111000100: data = 6'b111111;
12'b0010111000101: data = 6'b111111;
12'b0010111000110: data = 6'b111111;
12'b0010111000111: data = 6'b111111;
12'b0010111001000: data = 6'b111111;
12'b0010111001001: data = 6'b111111;
12'b0010111001010: data = 6'b111111;
12'b0010111001011: data = 6'b111111;
12'b0010111001100: data = 6'b111111;
12'b0010111001101: data = 6'b111111;
12'b0010111001110: data = 6'b111111;
12'b0010111001111: data = 6'b111111;
12'b0010111010000: data = 6'b111111;
12'b0010111010001: data = 6'b111111;
12'b0010111010010: data = 6'b111111;
12'b0010111010011: data = 6'b111111;
12'b0010111010100: data = 6'b111111;
12'b0010111010101: data = 6'b111111;
12'b0010111010110: data = 6'b111111;
12'b0010111010111: data = 6'b111111;
12'b0010111011000: data = 6'b111111;
12'b0010111011001: data = 6'b111111;
12'b0010111011010: data = 6'b111111;
12'b0010111011011: data = 6'b111111;
12'b0010111011100: data = 6'b111111;
12'b0010111011101: data = 6'b111111;
12'b0010111011110: data = 6'b111111;
12'b0010111011111: data = 6'b111111;
12'b0010111100000: data = 6'b111111;
12'b0010111100001: data = 6'b111111;
12'b0010111100010: data = 6'b111111;
12'b0010111100011: data = 6'b111111;
12'b0010111100100: data = 6'b111111;
12'b0010111100101: data = 6'b111111;
12'b0010111100110: data = 6'b111111;
12'b0010111100111: data = 6'b111111;
12'b0010111101000: data = 6'b111111;
12'b0010111101001: data = 6'b111111;
12'b0010111101010: data = 6'b111111;
12'b0010111101011: data = 6'b111111;
12'b0010111101100: data = 6'b111111;
12'b0010111101101: data = 6'b111111;
12'b0010111101110: data = 6'b111111;
12'b0010111101111: data = 6'b111111;
12'b0010111110000: data = 6'b111111;
12'b0010111110001: data = 6'b111111;
12'b0010111110010: data = 6'b111111;
12'b0010111110011: data = 6'b111111;
12'b0010111110100: data = 6'b111111;
12'b0010111110101: data = 6'b111111;
12'b0010111110110: data = 6'b111111;
12'b0010111110111: data = 6'b111111;
12'b0010111111000: data = 6'b111111;
12'b0010111111001: data = 6'b111111;
12'b0010111111010: data = 6'b111111;
12'b0010111111011: data = 6'b111111;
12'b0010111111100: data = 6'b111111;
12'b0010111111101: data = 6'b111111;
12'b0010111111110: data = 6'b111111;
12'b0010111111111: data = 6'b111111;
12'b00101110000000: data = 6'b111111;
12'b00101110000001: data = 6'b111111;
12'b00101110000010: data = 6'b111111;
12'b00101110000011: data = 6'b111111;
12'b00101110000100: data = 6'b111111;
12'b00101110000101: data = 6'b111111;
12'b00101110000110: data = 6'b111111;
12'b00101110000111: data = 6'b111111;
12'b00101110001000: data = 6'b111111;
12'b00101110001001: data = 6'b111111;
12'b00101110001010: data = 6'b111111;
12'b00101110001011: data = 6'b010101;
12'b00101110001100: data = 6'b000000;
12'b00101110001101: data = 6'b000000;
12'b00101110001110: data = 6'b101010;
12'b00101110001111: data = 6'b101010;
12'b00101110010000: data = 6'b101010;
12'b00101110010001: data = 6'b101010;
12'b00101110010010: data = 6'b010101;
12'b00101110010011: data = 6'b010101;
12'b00101110010100: data = 6'b010101;
12'b00101110010101: data = 6'b010101;
12'b00101110010110: data = 6'b010101;
12'b00101110010111: data = 6'b010101;
12'b00101110011000: data = 6'b010101;
12'b00101110011001: data = 6'b010101;
12'b00101110011010: data = 6'b010101;
12'b00101110011011: data = 6'b010101;
12'b00101110011100: data = 6'b010101;
12'b00101110011101: data = 6'b010101;
12'b00101110011110: data = 6'b010101;
12'b00101110011111: data = 6'b010101;
12'b00101110100000: data = 6'b010101;
12'b00101110100001: data = 6'b010101;
12'b00101110100010: data = 6'b010101;
12'b00101110100011: data = 6'b010101;
12'b00101110100100: data = 6'b010101;
12'b00101110100101: data = 6'b010101;
12'b00101110100110: data = 6'b010101;
12'b00101110100111: data = 6'b010101;
12'b00101110101000: data = 6'b010101;
12'b00101110101001: data = 6'b010101;
12'b00101110101010: data = 6'b010101;
12'b001100000000: data = 6'b010101;
12'b001100000001: data = 6'b010101;
12'b001100000010: data = 6'b010101;
12'b001100000011: data = 6'b010101;
12'b001100000100: data = 6'b010101;
12'b001100000101: data = 6'b010101;
12'b001100000110: data = 6'b010101;
12'b001100000111: data = 6'b010101;
12'b001100001000: data = 6'b010101;
12'b001100001001: data = 6'b010101;
12'b001100001010: data = 6'b010101;
12'b001100001011: data = 6'b010101;
12'b001100001100: data = 6'b010101;
12'b001100001101: data = 6'b010101;
12'b001100001110: data = 6'b010101;
12'b001100001111: data = 6'b010101;
12'b001100010000: data = 6'b010101;
12'b001100010001: data = 6'b010101;
12'b001100010010: data = 6'b010101;
12'b001100010011: data = 6'b010101;
12'b001100010100: data = 6'b010101;
12'b001100010101: data = 6'b010101;
12'b001100010110: data = 6'b010101;
12'b001100010111: data = 6'b010101;
12'b001100011000: data = 6'b010101;
12'b001100011001: data = 6'b101010;
12'b001100011010: data = 6'b101010;
12'b001100011011: data = 6'b101010;
12'b001100011100: data = 6'b010101;
12'b001100011101: data = 6'b000000;
12'b001100011110: data = 6'b000000;
12'b001100011111: data = 6'b010101;
12'b001100100000: data = 6'b111111;
12'b001100100001: data = 6'b111111;
12'b001100100010: data = 6'b111111;
12'b001100100011: data = 6'b111111;
12'b001100100100: data = 6'b111111;
12'b001100100101: data = 6'b111111;
12'b001100100110: data = 6'b111111;
12'b001100100111: data = 6'b111111;
12'b001100101000: data = 6'b111111;
12'b001100101001: data = 6'b111111;
12'b001100101010: data = 6'b111111;
12'b001100101011: data = 6'b111111;
12'b001100101100: data = 6'b111111;
12'b001100101101: data = 6'b111111;
12'b001100101110: data = 6'b111111;
12'b001100101111: data = 6'b111111;
12'b001100110000: data = 6'b111111;
12'b001100110001: data = 6'b111111;
12'b001100110010: data = 6'b111111;
12'b001100110011: data = 6'b111111;
12'b001100110100: data = 6'b111111;
12'b001100110101: data = 6'b111111;
12'b001100110110: data = 6'b111111;
12'b001100110111: data = 6'b111111;
12'b001100111000: data = 6'b111111;
12'b001100111001: data = 6'b111111;
12'b001100111010: data = 6'b111111;
12'b001100111011: data = 6'b111111;
12'b001100111100: data = 6'b111111;
12'b001100111101: data = 6'b111111;
12'b001100111110: data = 6'b111111;
12'b001100111111: data = 6'b111111;
12'b0011001000000: data = 6'b111111;
12'b0011001000001: data = 6'b111111;
12'b0011001000010: data = 6'b111111;
12'b0011001000011: data = 6'b111111;
12'b0011001000100: data = 6'b111111;
12'b0011001000101: data = 6'b111111;
12'b0011001000110: data = 6'b111111;
12'b0011001000111: data = 6'b111111;
12'b0011001001000: data = 6'b111111;
12'b0011001001001: data = 6'b111111;
12'b0011001001010: data = 6'b111111;
12'b0011001001011: data = 6'b111111;
12'b0011001001100: data = 6'b111111;
12'b0011001001101: data = 6'b111111;
12'b0011001001110: data = 6'b111111;
12'b0011001001111: data = 6'b111111;
12'b0011001010000: data = 6'b111111;
12'b0011001010001: data = 6'b111111;
12'b0011001010010: data = 6'b111111;
12'b0011001010011: data = 6'b111111;
12'b0011001010100: data = 6'b111111;
12'b0011001010101: data = 6'b111111;
12'b0011001010110: data = 6'b111111;
12'b0011001010111: data = 6'b111111;
12'b0011001011000: data = 6'b111111;
12'b0011001011001: data = 6'b111111;
12'b0011001011010: data = 6'b111111;
12'b0011001011011: data = 6'b111111;
12'b0011001011100: data = 6'b111111;
12'b0011001011101: data = 6'b111111;
12'b0011001011110: data = 6'b111111;
12'b0011001011111: data = 6'b111111;
12'b0011001100000: data = 6'b111111;
12'b0011001100001: data = 6'b111111;
12'b0011001100010: data = 6'b111111;
12'b0011001100011: data = 6'b111111;
12'b0011001100100: data = 6'b111111;
12'b0011001100101: data = 6'b111111;
12'b0011001100110: data = 6'b111111;
12'b0011001100111: data = 6'b111111;
12'b0011001101000: data = 6'b111111;
12'b0011001101001: data = 6'b111111;
12'b0011001101010: data = 6'b111111;
12'b0011001101011: data = 6'b111111;
12'b0011001101100: data = 6'b111111;
12'b0011001101101: data = 6'b111111;
12'b0011001101110: data = 6'b111111;
12'b0011001101111: data = 6'b111111;
12'b0011001110000: data = 6'b111111;
12'b0011001110001: data = 6'b111111;
12'b0011001110010: data = 6'b111111;
12'b0011001110011: data = 6'b111111;
12'b0011001110100: data = 6'b111111;
12'b0011001110101: data = 6'b111111;
12'b0011001110110: data = 6'b111111;
12'b0011001110111: data = 6'b111111;
12'b0011001111000: data = 6'b111111;
12'b0011001111001: data = 6'b111111;
12'b0011001111010: data = 6'b111111;
12'b0011001111011: data = 6'b111111;
12'b0011001111100: data = 6'b111111;
12'b0011001111101: data = 6'b111111;
12'b0011001111110: data = 6'b111111;
12'b0011001111111: data = 6'b111111;
12'b00110010000000: data = 6'b111111;
12'b00110010000001: data = 6'b111111;
12'b00110010000010: data = 6'b111111;
12'b00110010000011: data = 6'b111111;
12'b00110010000100: data = 6'b111111;
12'b00110010000101: data = 6'b111111;
12'b00110010000110: data = 6'b111111;
12'b00110010000111: data = 6'b111111;
12'b00110010001000: data = 6'b111111;
12'b00110010001001: data = 6'b111111;
12'b00110010001010: data = 6'b111111;
12'b00110010001011: data = 6'b010101;
12'b00110010001100: data = 6'b000000;
12'b00110010001101: data = 6'b000000;
12'b00110010001110: data = 6'b101010;
12'b00110010001111: data = 6'b101010;
12'b00110010010000: data = 6'b101010;
12'b00110010010001: data = 6'b101010;
12'b00110010010010: data = 6'b010101;
12'b00110010010011: data = 6'b010101;
12'b00110010010100: data = 6'b010101;
12'b00110010010101: data = 6'b010101;
12'b00110010010110: data = 6'b010101;
12'b00110010010111: data = 6'b010101;
12'b00110010011000: data = 6'b010101;
12'b00110010011001: data = 6'b010101;
12'b00110010011010: data = 6'b010101;
12'b00110010011011: data = 6'b010101;
12'b00110010011100: data = 6'b010101;
12'b00110010011101: data = 6'b010101;
12'b00110010011110: data = 6'b010101;
12'b00110010011111: data = 6'b010101;
12'b00110010100000: data = 6'b010101;
12'b00110010100001: data = 6'b010101;
12'b00110010100010: data = 6'b010101;
12'b00110010100011: data = 6'b010101;
12'b00110010100100: data = 6'b010101;
12'b00110010100101: data = 6'b010101;
12'b00110010100110: data = 6'b010101;
12'b00110010100111: data = 6'b010101;
12'b00110010101000: data = 6'b010101;
12'b00110010101001: data = 6'b010101;
12'b00110010101010: data = 6'b010101;
12'b001101000000: data = 6'b010101;
12'b001101000001: data = 6'b010101;
12'b001101000010: data = 6'b010101;
12'b001101000011: data = 6'b010101;
12'b001101000100: data = 6'b010101;
12'b001101000101: data = 6'b010101;
12'b001101000110: data = 6'b010101;
12'b001101000111: data = 6'b010101;
12'b001101001000: data = 6'b010101;
12'b001101001001: data = 6'b010101;
12'b001101001010: data = 6'b010101;
12'b001101001011: data = 6'b010101;
12'b001101001100: data = 6'b010101;
12'b001101001101: data = 6'b010101;
12'b001101001110: data = 6'b010101;
12'b001101001111: data = 6'b010101;
12'b001101010000: data = 6'b010101;
12'b001101010001: data = 6'b010101;
12'b001101010010: data = 6'b010101;
12'b001101010011: data = 6'b010101;
12'b001101010100: data = 6'b010101;
12'b001101010101: data = 6'b010101;
12'b001101010110: data = 6'b010101;
12'b001101010111: data = 6'b010101;
12'b001101011000: data = 6'b010101;
12'b001101011001: data = 6'b101010;
12'b001101011010: data = 6'b101010;
12'b001101011011: data = 6'b101010;
12'b001101011100: data = 6'b010101;
12'b001101011101: data = 6'b000000;
12'b001101011110: data = 6'b000000;
12'b001101011111: data = 6'b010101;
12'b001101100000: data = 6'b111111;
12'b001101100001: data = 6'b111111;
12'b001101100010: data = 6'b111111;
12'b001101100011: data = 6'b111111;
12'b001101100100: data = 6'b111111;
12'b001101100101: data = 6'b111111;
12'b001101100110: data = 6'b111111;
12'b001101100111: data = 6'b111111;
12'b001101101000: data = 6'b111111;
12'b001101101001: data = 6'b111111;
12'b001101101010: data = 6'b111111;
12'b001101101011: data = 6'b111111;
12'b001101101100: data = 6'b111111;
12'b001101101101: data = 6'b111111;
12'b001101101110: data = 6'b111111;
12'b001101101111: data = 6'b111111;
12'b001101110000: data = 6'b111111;
12'b001101110001: data = 6'b111111;
12'b001101110010: data = 6'b111111;
12'b001101110011: data = 6'b111111;
12'b001101110100: data = 6'b111111;
12'b001101110101: data = 6'b111111;
12'b001101110110: data = 6'b111111;
12'b001101110111: data = 6'b111111;
12'b001101111000: data = 6'b111111;
12'b001101111001: data = 6'b111111;
12'b001101111010: data = 6'b111111;
12'b001101111011: data = 6'b111111;
12'b001101111100: data = 6'b111111;
12'b001101111101: data = 6'b111111;
12'b001101111110: data = 6'b111111;
12'b001101111111: data = 6'b111111;
12'b0011011000000: data = 6'b111111;
12'b0011011000001: data = 6'b111111;
12'b0011011000010: data = 6'b111111;
12'b0011011000011: data = 6'b111111;
12'b0011011000100: data = 6'b111111;
12'b0011011000101: data = 6'b111111;
12'b0011011000110: data = 6'b111111;
12'b0011011000111: data = 6'b111111;
12'b0011011001000: data = 6'b111111;
12'b0011011001001: data = 6'b111111;
12'b0011011001010: data = 6'b111111;
12'b0011011001011: data = 6'b111111;
12'b0011011001100: data = 6'b111111;
12'b0011011001101: data = 6'b111111;
12'b0011011001110: data = 6'b111111;
12'b0011011001111: data = 6'b111111;
12'b0011011010000: data = 6'b111111;
12'b0011011010001: data = 6'b111111;
12'b0011011010010: data = 6'b111111;
12'b0011011010011: data = 6'b111111;
12'b0011011010100: data = 6'b111111;
12'b0011011010101: data = 6'b111111;
12'b0011011010110: data = 6'b111111;
12'b0011011010111: data = 6'b111111;
12'b0011011011000: data = 6'b111111;
12'b0011011011001: data = 6'b111111;
12'b0011011011010: data = 6'b111111;
12'b0011011011011: data = 6'b111111;
12'b0011011011100: data = 6'b111111;
12'b0011011011101: data = 6'b111111;
12'b0011011011110: data = 6'b111111;
12'b0011011011111: data = 6'b111111;
12'b0011011100000: data = 6'b111111;
12'b0011011100001: data = 6'b111111;
12'b0011011100010: data = 6'b111111;
12'b0011011100011: data = 6'b111111;
12'b0011011100100: data = 6'b111111;
12'b0011011100101: data = 6'b111111;
12'b0011011100110: data = 6'b111111;
12'b0011011100111: data = 6'b111111;
12'b0011011101000: data = 6'b111111;
12'b0011011101001: data = 6'b111111;
12'b0011011101010: data = 6'b111111;
12'b0011011101011: data = 6'b111111;
12'b0011011101100: data = 6'b111111;
12'b0011011101101: data = 6'b111111;
12'b0011011101110: data = 6'b111111;
12'b0011011101111: data = 6'b111111;
12'b0011011110000: data = 6'b111111;
12'b0011011110001: data = 6'b111111;
12'b0011011110010: data = 6'b111111;
12'b0011011110011: data = 6'b111111;
12'b0011011110100: data = 6'b111111;
12'b0011011110101: data = 6'b111111;
12'b0011011110110: data = 6'b111111;
12'b0011011110111: data = 6'b111111;
12'b0011011111000: data = 6'b111111;
12'b0011011111001: data = 6'b111111;
12'b0011011111010: data = 6'b111111;
12'b0011011111011: data = 6'b111111;
12'b0011011111100: data = 6'b111111;
12'b0011011111101: data = 6'b111111;
12'b0011011111110: data = 6'b111111;
12'b0011011111111: data = 6'b111111;
12'b00110110000000: data = 6'b111111;
12'b00110110000001: data = 6'b111111;
12'b00110110000010: data = 6'b111111;
12'b00110110000011: data = 6'b111111;
12'b00110110000100: data = 6'b111111;
12'b00110110000101: data = 6'b111111;
12'b00110110000110: data = 6'b111111;
12'b00110110000111: data = 6'b111111;
12'b00110110001000: data = 6'b111111;
12'b00110110001001: data = 6'b111111;
12'b00110110001010: data = 6'b111111;
12'b00110110001011: data = 6'b010101;
12'b00110110001100: data = 6'b000000;
12'b00110110001101: data = 6'b000000;
12'b00110110001110: data = 6'b101010;
12'b00110110001111: data = 6'b101010;
12'b00110110010000: data = 6'b101010;
12'b00110110010001: data = 6'b101010;
12'b00110110010010: data = 6'b010101;
12'b00110110010011: data = 6'b010101;
12'b00110110010100: data = 6'b010101;
12'b00110110010101: data = 6'b010101;
12'b00110110010110: data = 6'b010101;
12'b00110110010111: data = 6'b010101;
12'b00110110011000: data = 6'b010101;
12'b00110110011001: data = 6'b010101;
12'b00110110011010: data = 6'b010101;
12'b00110110011011: data = 6'b010101;
12'b00110110011100: data = 6'b010101;
12'b00110110011101: data = 6'b010101;
12'b00110110011110: data = 6'b010101;
12'b00110110011111: data = 6'b010101;
12'b00110110100000: data = 6'b010101;
12'b00110110100001: data = 6'b010101;
12'b00110110100010: data = 6'b010101;
12'b00110110100011: data = 6'b010101;
12'b00110110100100: data = 6'b010101;
12'b00110110100101: data = 6'b010101;
12'b00110110100110: data = 6'b010101;
12'b00110110100111: data = 6'b010101;
12'b00110110101000: data = 6'b010101;
12'b00110110101001: data = 6'b010101;
12'b00110110101010: data = 6'b010101;
12'b001110000000: data = 6'b010101;
12'b001110000001: data = 6'b010101;
12'b001110000010: data = 6'b010101;
12'b001110000011: data = 6'b010101;
12'b001110000100: data = 6'b010101;
12'b001110000101: data = 6'b010101;
12'b001110000110: data = 6'b010101;
12'b001110000111: data = 6'b010101;
12'b001110001000: data = 6'b010101;
12'b001110001001: data = 6'b010101;
12'b001110001010: data = 6'b010101;
12'b001110001011: data = 6'b010101;
12'b001110001100: data = 6'b010101;
12'b001110001101: data = 6'b010101;
12'b001110001110: data = 6'b010101;
12'b001110001111: data = 6'b010101;
12'b001110010000: data = 6'b010101;
12'b001110010001: data = 6'b010101;
12'b001110010010: data = 6'b010101;
12'b001110010011: data = 6'b010101;
12'b001110010100: data = 6'b010101;
12'b001110010101: data = 6'b010101;
12'b001110010110: data = 6'b010101;
12'b001110010111: data = 6'b010101;
12'b001110011000: data = 6'b010101;
12'b001110011001: data = 6'b101010;
12'b001110011010: data = 6'b101010;
12'b001110011011: data = 6'b101010;
12'b001110011100: data = 6'b010101;
12'b001110011101: data = 6'b000000;
12'b001110011110: data = 6'b000000;
12'b001110011111: data = 6'b010101;
12'b001110100000: data = 6'b111111;
12'b001110100001: data = 6'b111111;
12'b001110100010: data = 6'b111111;
12'b001110100011: data = 6'b111111;
12'b001110100100: data = 6'b111111;
12'b001110100101: data = 6'b111111;
12'b001110100110: data = 6'b111111;
12'b001110100111: data = 6'b111111;
12'b001110101000: data = 6'b111111;
12'b001110101001: data = 6'b111111;
12'b001110101010: data = 6'b111111;
12'b001110101011: data = 6'b111111;
12'b001110101100: data = 6'b111111;
12'b001110101101: data = 6'b111111;
12'b001110101110: data = 6'b111111;
12'b001110101111: data = 6'b111111;
12'b001110110000: data = 6'b111111;
12'b001110110001: data = 6'b111111;
12'b001110110010: data = 6'b111111;
12'b001110110011: data = 6'b111111;
12'b001110110100: data = 6'b111111;
12'b001110110101: data = 6'b111111;
12'b001110110110: data = 6'b111111;
12'b001110110111: data = 6'b111111;
12'b001110111000: data = 6'b111111;
12'b001110111001: data = 6'b111111;
12'b001110111010: data = 6'b111111;
12'b001110111011: data = 6'b111111;
12'b001110111100: data = 6'b111111;
12'b001110111101: data = 6'b111111;
12'b001110111110: data = 6'b111111;
12'b001110111111: data = 6'b111111;
12'b0011101000000: data = 6'b111111;
12'b0011101000001: data = 6'b111111;
12'b0011101000010: data = 6'b111111;
12'b0011101000011: data = 6'b111111;
12'b0011101000100: data = 6'b111111;
12'b0011101000101: data = 6'b111111;
12'b0011101000110: data = 6'b111111;
12'b0011101000111: data = 6'b111111;
12'b0011101001000: data = 6'b111111;
12'b0011101001001: data = 6'b111111;
12'b0011101001010: data = 6'b111111;
12'b0011101001011: data = 6'b111111;
12'b0011101001100: data = 6'b111111;
12'b0011101001101: data = 6'b111111;
12'b0011101001110: data = 6'b111111;
12'b0011101001111: data = 6'b111111;
12'b0011101010000: data = 6'b111111;
12'b0011101010001: data = 6'b111111;
12'b0011101010010: data = 6'b111111;
12'b0011101010011: data = 6'b111111;
12'b0011101010100: data = 6'b111111;
12'b0011101010101: data = 6'b111111;
12'b0011101010110: data = 6'b111111;
12'b0011101010111: data = 6'b111111;
12'b0011101011000: data = 6'b111111;
12'b0011101011001: data = 6'b111111;
12'b0011101011010: data = 6'b111111;
12'b0011101011011: data = 6'b111111;
12'b0011101011100: data = 6'b111111;
12'b0011101011101: data = 6'b111111;
12'b0011101011110: data = 6'b111111;
12'b0011101011111: data = 6'b111111;
12'b0011101100000: data = 6'b111111;
12'b0011101100001: data = 6'b111111;
12'b0011101100010: data = 6'b111111;
12'b0011101100011: data = 6'b111111;
12'b0011101100100: data = 6'b111111;
12'b0011101100101: data = 6'b111111;
12'b0011101100110: data = 6'b111111;
12'b0011101100111: data = 6'b111111;
12'b0011101101000: data = 6'b111111;
12'b0011101101001: data = 6'b111111;
12'b0011101101010: data = 6'b111111;
12'b0011101101011: data = 6'b111111;
12'b0011101101100: data = 6'b111111;
12'b0011101101101: data = 6'b111111;
12'b0011101101110: data = 6'b111111;
12'b0011101101111: data = 6'b111111;
12'b0011101110000: data = 6'b111111;
12'b0011101110001: data = 6'b111111;
12'b0011101110010: data = 6'b111111;
12'b0011101110011: data = 6'b111111;
12'b0011101110100: data = 6'b111111;
12'b0011101110101: data = 6'b111111;
12'b0011101110110: data = 6'b111111;
12'b0011101110111: data = 6'b111111;
12'b0011101111000: data = 6'b111111;
12'b0011101111001: data = 6'b111111;
12'b0011101111010: data = 6'b111111;
12'b0011101111011: data = 6'b111111;
12'b0011101111100: data = 6'b111111;
12'b0011101111101: data = 6'b111111;
12'b0011101111110: data = 6'b111111;
12'b0011101111111: data = 6'b111111;
12'b00111010000000: data = 6'b111111;
12'b00111010000001: data = 6'b111111;
12'b00111010000010: data = 6'b111111;
12'b00111010000011: data = 6'b111111;
12'b00111010000100: data = 6'b111111;
12'b00111010000101: data = 6'b111111;
12'b00111010000110: data = 6'b111111;
12'b00111010000111: data = 6'b111111;
12'b00111010001000: data = 6'b111111;
12'b00111010001001: data = 6'b111111;
12'b00111010001010: data = 6'b111111;
12'b00111010001011: data = 6'b010101;
12'b00111010001100: data = 6'b000000;
12'b00111010001101: data = 6'b000000;
12'b00111010001110: data = 6'b101010;
12'b00111010001111: data = 6'b101010;
12'b00111010010000: data = 6'b101010;
12'b00111010010001: data = 6'b101010;
12'b00111010010010: data = 6'b010101;
12'b00111010010011: data = 6'b010101;
12'b00111010010100: data = 6'b010101;
12'b00111010010101: data = 6'b010101;
12'b00111010010110: data = 6'b010101;
12'b00111010010111: data = 6'b010101;
12'b00111010011000: data = 6'b010101;
12'b00111010011001: data = 6'b010101;
12'b00111010011010: data = 6'b010101;
12'b00111010011011: data = 6'b010101;
12'b00111010011100: data = 6'b010101;
12'b00111010011101: data = 6'b010101;
12'b00111010011110: data = 6'b010101;
12'b00111010011111: data = 6'b010101;
12'b00111010100000: data = 6'b010101;
12'b00111010100001: data = 6'b010101;
12'b00111010100010: data = 6'b010101;
12'b00111010100011: data = 6'b010101;
12'b00111010100100: data = 6'b010101;
12'b00111010100101: data = 6'b010101;
12'b00111010100110: data = 6'b010101;
12'b00111010100111: data = 6'b010101;
12'b00111010101000: data = 6'b010101;
12'b00111010101001: data = 6'b010101;
12'b00111010101010: data = 6'b010101;
12'b001111000000: data = 6'b010101;
12'b001111000001: data = 6'b010101;
12'b001111000010: data = 6'b010101;
12'b001111000011: data = 6'b010101;
12'b001111000100: data = 6'b010101;
12'b001111000101: data = 6'b010101;
12'b001111000110: data = 6'b010101;
12'b001111000111: data = 6'b010101;
12'b001111001000: data = 6'b010101;
12'b001111001001: data = 6'b010101;
12'b001111001010: data = 6'b010101;
12'b001111001011: data = 6'b010101;
12'b001111001100: data = 6'b010101;
12'b001111001101: data = 6'b010101;
12'b001111001110: data = 6'b010101;
12'b001111001111: data = 6'b010101;
12'b001111010000: data = 6'b010101;
12'b001111010001: data = 6'b010101;
12'b001111010010: data = 6'b010101;
12'b001111010011: data = 6'b010101;
12'b001111010100: data = 6'b010101;
12'b001111010101: data = 6'b010101;
12'b001111010110: data = 6'b010101;
12'b001111010111: data = 6'b010101;
12'b001111011000: data = 6'b010101;
12'b001111011001: data = 6'b101010;
12'b001111011010: data = 6'b101010;
12'b001111011011: data = 6'b101010;
12'b001111011100: data = 6'b010101;
12'b001111011101: data = 6'b000000;
12'b001111011110: data = 6'b000000;
12'b001111011111: data = 6'b010101;
12'b001111100000: data = 6'b111111;
12'b001111100001: data = 6'b111111;
12'b001111100010: data = 6'b111111;
12'b001111100011: data = 6'b111111;
12'b001111100100: data = 6'b111111;
12'b001111100101: data = 6'b111111;
12'b001111100110: data = 6'b111111;
12'b001111100111: data = 6'b111111;
12'b001111101000: data = 6'b111111;
12'b001111101001: data = 6'b111111;
12'b001111101010: data = 6'b111111;
12'b001111101011: data = 6'b111111;
12'b001111101100: data = 6'b111111;
12'b001111101101: data = 6'b111111;
12'b001111101110: data = 6'b111111;
12'b001111101111: data = 6'b111111;
12'b001111110000: data = 6'b111111;
12'b001111110001: data = 6'b111111;
12'b001111110010: data = 6'b111111;
12'b001111110011: data = 6'b111111;
12'b001111110100: data = 6'b111111;
12'b001111110101: data = 6'b111111;
12'b001111110110: data = 6'b111111;
12'b001111110111: data = 6'b111111;
12'b001111111000: data = 6'b111111;
12'b001111111001: data = 6'b111111;
12'b001111111010: data = 6'b111111;
12'b001111111011: data = 6'b111111;
12'b001111111100: data = 6'b111111;
12'b001111111101: data = 6'b111111;
12'b001111111110: data = 6'b111111;
12'b001111111111: data = 6'b111111;
12'b0011111000000: data = 6'b111111;
12'b0011111000001: data = 6'b111111;
12'b0011111000010: data = 6'b111111;
12'b0011111000011: data = 6'b111111;
12'b0011111000100: data = 6'b111111;
12'b0011111000101: data = 6'b111111;
12'b0011111000110: data = 6'b111111;
12'b0011111000111: data = 6'b111111;
12'b0011111001000: data = 6'b111111;
12'b0011111001001: data = 6'b111111;
12'b0011111001010: data = 6'b111111;
12'b0011111001011: data = 6'b111111;
12'b0011111001100: data = 6'b111111;
12'b0011111001101: data = 6'b111111;
12'b0011111001110: data = 6'b111111;
12'b0011111001111: data = 6'b111111;
12'b0011111010000: data = 6'b111111;
12'b0011111010001: data = 6'b111111;
12'b0011111010010: data = 6'b111111;
12'b0011111010011: data = 6'b111111;
12'b0011111010100: data = 6'b111111;
12'b0011111010101: data = 6'b111111;
12'b0011111010110: data = 6'b111111;
12'b0011111010111: data = 6'b111111;
12'b0011111011000: data = 6'b111111;
12'b0011111011001: data = 6'b111111;
12'b0011111011010: data = 6'b111111;
12'b0011111011011: data = 6'b111111;
12'b0011111011100: data = 6'b111111;
12'b0011111011101: data = 6'b111111;
12'b0011111011110: data = 6'b111111;
12'b0011111011111: data = 6'b111111;
12'b0011111100000: data = 6'b111111;
12'b0011111100001: data = 6'b111111;
12'b0011111100010: data = 6'b111111;
12'b0011111100011: data = 6'b111111;
12'b0011111100100: data = 6'b111111;
12'b0011111100101: data = 6'b111111;
12'b0011111100110: data = 6'b111111;
12'b0011111100111: data = 6'b111111;
12'b0011111101000: data = 6'b111111;
12'b0011111101001: data = 6'b111111;
12'b0011111101010: data = 6'b111111;
12'b0011111101011: data = 6'b111111;
12'b0011111101100: data = 6'b111111;
12'b0011111101101: data = 6'b111111;
12'b0011111101110: data = 6'b111111;
12'b0011111101111: data = 6'b111111;
12'b0011111110000: data = 6'b111111;
12'b0011111110001: data = 6'b111111;
12'b0011111110010: data = 6'b111111;
12'b0011111110011: data = 6'b111111;
12'b0011111110100: data = 6'b111111;
12'b0011111110101: data = 6'b111111;
12'b0011111110110: data = 6'b111111;
12'b0011111110111: data = 6'b111111;
12'b0011111111000: data = 6'b111111;
12'b0011111111001: data = 6'b111111;
12'b0011111111010: data = 6'b111111;
12'b0011111111011: data = 6'b111111;
12'b0011111111100: data = 6'b111111;
12'b0011111111101: data = 6'b111111;
12'b0011111111110: data = 6'b111111;
12'b0011111111111: data = 6'b111111;
12'b00111110000000: data = 6'b111111;
12'b00111110000001: data = 6'b111111;
12'b00111110000010: data = 6'b111111;
12'b00111110000011: data = 6'b111111;
12'b00111110000100: data = 6'b111111;
12'b00111110000101: data = 6'b111111;
12'b00111110000110: data = 6'b111111;
12'b00111110000111: data = 6'b111111;
12'b00111110001000: data = 6'b111111;
12'b00111110001001: data = 6'b111111;
12'b00111110001010: data = 6'b111111;
12'b00111110001011: data = 6'b010101;
12'b00111110001100: data = 6'b000000;
12'b00111110001101: data = 6'b000000;
12'b00111110001110: data = 6'b101010;
12'b00111110001111: data = 6'b101010;
12'b00111110010000: data = 6'b101010;
12'b00111110010001: data = 6'b101010;
12'b00111110010010: data = 6'b010101;
12'b00111110010011: data = 6'b010101;
12'b00111110010100: data = 6'b010101;
12'b00111110010101: data = 6'b010101;
12'b00111110010110: data = 6'b010101;
12'b00111110010111: data = 6'b010101;
12'b00111110011000: data = 6'b010101;
12'b00111110011001: data = 6'b010101;
12'b00111110011010: data = 6'b010101;
12'b00111110011011: data = 6'b010101;
12'b00111110011100: data = 6'b010101;
12'b00111110011101: data = 6'b010101;
12'b00111110011110: data = 6'b010101;
12'b00111110011111: data = 6'b010101;
12'b00111110100000: data = 6'b010101;
12'b00111110100001: data = 6'b010101;
12'b00111110100010: data = 6'b010101;
12'b00111110100011: data = 6'b010101;
12'b00111110100100: data = 6'b010101;
12'b00111110100101: data = 6'b010101;
12'b00111110100110: data = 6'b010101;
12'b00111110100111: data = 6'b010101;
12'b00111110101000: data = 6'b010101;
12'b00111110101001: data = 6'b010101;
12'b00111110101010: data = 6'b010101;
12'b010000000000: data = 6'b010101;
12'b010000000001: data = 6'b010101;
12'b010000000010: data = 6'b010101;
12'b010000000011: data = 6'b010101;
12'b010000000100: data = 6'b010101;
12'b010000000101: data = 6'b010101;
12'b010000000110: data = 6'b010101;
12'b010000000111: data = 6'b010101;
12'b010000001000: data = 6'b010101;
12'b010000001001: data = 6'b010101;
12'b010000001010: data = 6'b010101;
12'b010000001011: data = 6'b010101;
12'b010000001100: data = 6'b010101;
12'b010000001101: data = 6'b010101;
12'b010000001110: data = 6'b010101;
12'b010000001111: data = 6'b010101;
12'b010000010000: data = 6'b010101;
12'b010000010001: data = 6'b010101;
12'b010000010010: data = 6'b010101;
12'b010000010011: data = 6'b010101;
12'b010000010100: data = 6'b010101;
12'b010000010101: data = 6'b010101;
12'b010000010110: data = 6'b010101;
12'b010000010111: data = 6'b010101;
12'b010000011000: data = 6'b010101;
12'b010000011001: data = 6'b101010;
12'b010000011010: data = 6'b101010;
12'b010000011011: data = 6'b101010;
12'b010000011100: data = 6'b010101;
12'b010000011101: data = 6'b000000;
12'b010000011110: data = 6'b000000;
12'b010000011111: data = 6'b010101;
12'b010000100000: data = 6'b111111;
12'b010000100001: data = 6'b111111;
12'b010000100010: data = 6'b111111;
12'b010000100011: data = 6'b111111;
12'b010000100100: data = 6'b111111;
12'b010000100101: data = 6'b111111;
12'b010000100110: data = 6'b111111;
12'b010000100111: data = 6'b111111;
12'b010000101000: data = 6'b111111;
12'b010000101001: data = 6'b111111;
12'b010000101010: data = 6'b111111;
12'b010000101011: data = 6'b111111;
12'b010000101100: data = 6'b111111;
12'b010000101101: data = 6'b111111;
12'b010000101110: data = 6'b111111;
12'b010000101111: data = 6'b111111;
12'b010000110000: data = 6'b111111;
12'b010000110001: data = 6'b111111;
12'b010000110010: data = 6'b111111;
12'b010000110011: data = 6'b111111;
12'b010000110100: data = 6'b111111;
12'b010000110101: data = 6'b111111;
12'b010000110110: data = 6'b111111;
12'b010000110111: data = 6'b111111;
12'b010000111000: data = 6'b111111;
12'b010000111001: data = 6'b111111;
12'b010000111010: data = 6'b111111;
12'b010000111011: data = 6'b111111;
12'b010000111100: data = 6'b111111;
12'b010000111101: data = 6'b111111;
12'b010000111110: data = 6'b111111;
12'b010000111111: data = 6'b111111;
12'b0100001000000: data = 6'b111111;
12'b0100001000001: data = 6'b111111;
12'b0100001000010: data = 6'b111111;
12'b0100001000011: data = 6'b111111;
12'b0100001000100: data = 6'b111111;
12'b0100001000101: data = 6'b111111;
12'b0100001000110: data = 6'b111111;
12'b0100001000111: data = 6'b111111;
12'b0100001001000: data = 6'b111111;
12'b0100001001001: data = 6'b111111;
12'b0100001001010: data = 6'b111111;
12'b0100001001011: data = 6'b111111;
12'b0100001001100: data = 6'b111111;
12'b0100001001101: data = 6'b111111;
12'b0100001001110: data = 6'b111111;
12'b0100001001111: data = 6'b111111;
12'b0100001010000: data = 6'b111111;
12'b0100001010001: data = 6'b111111;
12'b0100001010010: data = 6'b111111;
12'b0100001010011: data = 6'b111111;
12'b0100001010100: data = 6'b111111;
12'b0100001010101: data = 6'b111111;
12'b0100001010110: data = 6'b111111;
12'b0100001010111: data = 6'b111111;
12'b0100001011000: data = 6'b111111;
12'b0100001011001: data = 6'b111111;
12'b0100001011010: data = 6'b111111;
12'b0100001011011: data = 6'b111111;
12'b0100001011100: data = 6'b111111;
12'b0100001011101: data = 6'b111111;
12'b0100001011110: data = 6'b111111;
12'b0100001011111: data = 6'b111111;
12'b0100001100000: data = 6'b111111;
12'b0100001100001: data = 6'b111111;
12'b0100001100010: data = 6'b111111;
12'b0100001100011: data = 6'b111111;
12'b0100001100100: data = 6'b111111;
12'b0100001100101: data = 6'b111111;
12'b0100001100110: data = 6'b111111;
12'b0100001100111: data = 6'b111111;
12'b0100001101000: data = 6'b111111;
12'b0100001101001: data = 6'b111111;
12'b0100001101010: data = 6'b111111;
12'b0100001101011: data = 6'b111111;
12'b0100001101100: data = 6'b111111;
12'b0100001101101: data = 6'b111111;
12'b0100001101110: data = 6'b111111;
12'b0100001101111: data = 6'b111111;
12'b0100001110000: data = 6'b111111;
12'b0100001110001: data = 6'b111111;
12'b0100001110010: data = 6'b111111;
12'b0100001110011: data = 6'b111111;
12'b0100001110100: data = 6'b111111;
12'b0100001110101: data = 6'b111111;
12'b0100001110110: data = 6'b111111;
12'b0100001110111: data = 6'b111111;
12'b0100001111000: data = 6'b111111;
12'b0100001111001: data = 6'b111111;
12'b0100001111010: data = 6'b111111;
12'b0100001111011: data = 6'b111111;
12'b0100001111100: data = 6'b111111;
12'b0100001111101: data = 6'b111111;
12'b0100001111110: data = 6'b111111;
12'b0100001111111: data = 6'b111111;
12'b01000010000000: data = 6'b111111;
12'b01000010000001: data = 6'b111111;
12'b01000010000010: data = 6'b111111;
12'b01000010000011: data = 6'b111111;
12'b01000010000100: data = 6'b111111;
12'b01000010000101: data = 6'b111111;
12'b01000010000110: data = 6'b111111;
12'b01000010000111: data = 6'b111111;
12'b01000010001000: data = 6'b111111;
12'b01000010001001: data = 6'b111111;
12'b01000010001010: data = 6'b111111;
12'b01000010001011: data = 6'b010101;
12'b01000010001100: data = 6'b000000;
12'b01000010001101: data = 6'b000000;
12'b01000010001110: data = 6'b101010;
12'b01000010001111: data = 6'b101010;
12'b01000010010000: data = 6'b101010;
12'b01000010010001: data = 6'b101010;
12'b01000010010010: data = 6'b010101;
12'b01000010010011: data = 6'b010101;
12'b01000010010100: data = 6'b010101;
12'b01000010010101: data = 6'b010101;
12'b01000010010110: data = 6'b010101;
12'b01000010010111: data = 6'b010101;
12'b01000010011000: data = 6'b010101;
12'b01000010011001: data = 6'b010101;
12'b01000010011010: data = 6'b010101;
12'b01000010011011: data = 6'b010101;
12'b01000010011100: data = 6'b010101;
12'b01000010011101: data = 6'b010101;
12'b01000010011110: data = 6'b010101;
12'b01000010011111: data = 6'b010101;
12'b01000010100000: data = 6'b010101;
12'b01000010100001: data = 6'b010101;
12'b01000010100010: data = 6'b010101;
12'b01000010100011: data = 6'b010101;
12'b01000010100100: data = 6'b010101;
12'b01000010100101: data = 6'b010101;
12'b01000010100110: data = 6'b010101;
12'b01000010100111: data = 6'b010101;
12'b01000010101000: data = 6'b010101;
12'b01000010101001: data = 6'b010101;
12'b01000010101010: data = 6'b010101;
12'b010001000000: data = 6'b010101;
12'b010001000001: data = 6'b010101;
12'b010001000010: data = 6'b010101;
12'b010001000011: data = 6'b010101;
12'b010001000100: data = 6'b010101;
12'b010001000101: data = 6'b010101;
12'b010001000110: data = 6'b010101;
12'b010001000111: data = 6'b010101;
12'b010001001000: data = 6'b010101;
12'b010001001001: data = 6'b010101;
12'b010001001010: data = 6'b010101;
12'b010001001011: data = 6'b010101;
12'b010001001100: data = 6'b010101;
12'b010001001101: data = 6'b010101;
12'b010001001110: data = 6'b010101;
12'b010001001111: data = 6'b010101;
12'b010001010000: data = 6'b010101;
12'b010001010001: data = 6'b010101;
12'b010001010010: data = 6'b010101;
12'b010001010011: data = 6'b010101;
12'b010001010100: data = 6'b010101;
12'b010001010101: data = 6'b010101;
12'b010001010110: data = 6'b010101;
12'b010001010111: data = 6'b010101;
12'b010001011000: data = 6'b010101;
12'b010001011001: data = 6'b101010;
12'b010001011010: data = 6'b101010;
12'b010001011011: data = 6'b101010;
12'b010001011100: data = 6'b010101;
12'b010001011101: data = 6'b000000;
12'b010001011110: data = 6'b000000;
12'b010001011111: data = 6'b010101;
12'b010001100000: data = 6'b111111;
12'b010001100001: data = 6'b111111;
12'b010001100010: data = 6'b111111;
12'b010001100011: data = 6'b111111;
12'b010001100100: data = 6'b111111;
12'b010001100101: data = 6'b111111;
12'b010001100110: data = 6'b111111;
12'b010001100111: data = 6'b111111;
12'b010001101000: data = 6'b111111;
12'b010001101001: data = 6'b111111;
12'b010001101010: data = 6'b111111;
12'b010001101011: data = 6'b111111;
12'b010001101100: data = 6'b111111;
12'b010001101101: data = 6'b111111;
12'b010001101110: data = 6'b111111;
12'b010001101111: data = 6'b111111;
12'b010001110000: data = 6'b111111;
12'b010001110001: data = 6'b111111;
12'b010001110010: data = 6'b111111;
12'b010001110011: data = 6'b111111;
12'b010001110100: data = 6'b111111;
12'b010001110101: data = 6'b111111;
12'b010001110110: data = 6'b111111;
12'b010001110111: data = 6'b111111;
12'b010001111000: data = 6'b111111;
12'b010001111001: data = 6'b111111;
12'b010001111010: data = 6'b111111;
12'b010001111011: data = 6'b111111;
12'b010001111100: data = 6'b111111;
12'b010001111101: data = 6'b111111;
12'b010001111110: data = 6'b111111;
12'b010001111111: data = 6'b111111;
12'b0100011000000: data = 6'b111111;
12'b0100011000001: data = 6'b111111;
12'b0100011000010: data = 6'b111111;
12'b0100011000011: data = 6'b111111;
12'b0100011000100: data = 6'b111111;
12'b0100011000101: data = 6'b111111;
12'b0100011000110: data = 6'b111111;
12'b0100011000111: data = 6'b111111;
12'b0100011001000: data = 6'b111111;
12'b0100011001001: data = 6'b111111;
12'b0100011001010: data = 6'b111111;
12'b0100011001011: data = 6'b111111;
12'b0100011001100: data = 6'b111111;
12'b0100011001101: data = 6'b111111;
12'b0100011001110: data = 6'b111111;
12'b0100011001111: data = 6'b111111;
12'b0100011010000: data = 6'b111111;
12'b0100011010001: data = 6'b111111;
12'b0100011010010: data = 6'b111111;
12'b0100011010011: data = 6'b111111;
12'b0100011010100: data = 6'b111111;
12'b0100011010101: data = 6'b111111;
12'b0100011010110: data = 6'b111111;
12'b0100011010111: data = 6'b111111;
12'b0100011011000: data = 6'b111111;
12'b0100011011001: data = 6'b111111;
12'b0100011011010: data = 6'b111111;
12'b0100011011011: data = 6'b111111;
12'b0100011011100: data = 6'b111111;
12'b0100011011101: data = 6'b111111;
12'b0100011011110: data = 6'b111111;
12'b0100011011111: data = 6'b111111;
12'b0100011100000: data = 6'b111111;
12'b0100011100001: data = 6'b111111;
12'b0100011100010: data = 6'b111111;
12'b0100011100011: data = 6'b111111;
12'b0100011100100: data = 6'b111111;
12'b0100011100101: data = 6'b111111;
12'b0100011100110: data = 6'b111111;
12'b0100011100111: data = 6'b111111;
12'b0100011101000: data = 6'b111111;
12'b0100011101001: data = 6'b111111;
12'b0100011101010: data = 6'b111111;
12'b0100011101011: data = 6'b111111;
12'b0100011101100: data = 6'b111111;
12'b0100011101101: data = 6'b111111;
12'b0100011101110: data = 6'b111111;
12'b0100011101111: data = 6'b111111;
12'b0100011110000: data = 6'b111111;
12'b0100011110001: data = 6'b111111;
12'b0100011110010: data = 6'b111111;
12'b0100011110011: data = 6'b111111;
12'b0100011110100: data = 6'b111111;
12'b0100011110101: data = 6'b111111;
12'b0100011110110: data = 6'b111111;
12'b0100011110111: data = 6'b111111;
12'b0100011111000: data = 6'b111111;
12'b0100011111001: data = 6'b111111;
12'b0100011111010: data = 6'b111111;
12'b0100011111011: data = 6'b111111;
12'b0100011111100: data = 6'b111111;
12'b0100011111101: data = 6'b111111;
12'b0100011111110: data = 6'b111111;
12'b0100011111111: data = 6'b111111;
12'b01000110000000: data = 6'b111111;
12'b01000110000001: data = 6'b111111;
12'b01000110000010: data = 6'b111111;
12'b01000110000011: data = 6'b111111;
12'b01000110000100: data = 6'b111111;
12'b01000110000101: data = 6'b111111;
12'b01000110000110: data = 6'b111111;
12'b01000110000111: data = 6'b111111;
12'b01000110001000: data = 6'b111111;
12'b01000110001001: data = 6'b111111;
12'b01000110001010: data = 6'b111111;
12'b01000110001011: data = 6'b010101;
12'b01000110001100: data = 6'b000000;
12'b01000110001101: data = 6'b000000;
12'b01000110001110: data = 6'b101010;
12'b01000110001111: data = 6'b101010;
12'b01000110010000: data = 6'b101010;
12'b01000110010001: data = 6'b101010;
12'b01000110010010: data = 6'b010101;
12'b01000110010011: data = 6'b010101;
12'b01000110010100: data = 6'b010101;
12'b01000110010101: data = 6'b010101;
12'b01000110010110: data = 6'b010101;
12'b01000110010111: data = 6'b010101;
12'b01000110011000: data = 6'b010101;
12'b01000110011001: data = 6'b010101;
12'b01000110011010: data = 6'b010101;
12'b01000110011011: data = 6'b010101;
12'b01000110011100: data = 6'b010101;
12'b01000110011101: data = 6'b010101;
12'b01000110011110: data = 6'b010101;
12'b01000110011111: data = 6'b010101;
12'b01000110100000: data = 6'b010101;
12'b01000110100001: data = 6'b010101;
12'b01000110100010: data = 6'b010101;
12'b01000110100011: data = 6'b010101;
12'b01000110100100: data = 6'b010101;
12'b01000110100101: data = 6'b010101;
12'b01000110100110: data = 6'b010101;
12'b01000110100111: data = 6'b010101;
12'b01000110101000: data = 6'b010101;
12'b01000110101001: data = 6'b010101;
12'b01000110101010: data = 6'b010101;
12'b010010000000: data = 6'b010101;
12'b010010000001: data = 6'b010101;
12'b010010000010: data = 6'b010101;
12'b010010000011: data = 6'b010101;
12'b010010000100: data = 6'b010101;
12'b010010000101: data = 6'b010101;
12'b010010000110: data = 6'b010101;
12'b010010000111: data = 6'b010101;
12'b010010001000: data = 6'b010101;
12'b010010001001: data = 6'b010101;
12'b010010001010: data = 6'b010101;
12'b010010001011: data = 6'b010101;
12'b010010001100: data = 6'b010101;
12'b010010001101: data = 6'b010101;
12'b010010001110: data = 6'b010101;
12'b010010001111: data = 6'b010101;
12'b010010010000: data = 6'b010101;
12'b010010010001: data = 6'b010101;
12'b010010010010: data = 6'b010101;
12'b010010010011: data = 6'b010101;
12'b010010010100: data = 6'b010101;
12'b010010010101: data = 6'b010101;
12'b010010010110: data = 6'b010101;
12'b010010010111: data = 6'b010101;
12'b010010011000: data = 6'b010101;
12'b010010011001: data = 6'b101010;
12'b010010011010: data = 6'b101010;
12'b010010011011: data = 6'b101010;
12'b010010011100: data = 6'b010101;
12'b010010011101: data = 6'b000000;
12'b010010011110: data = 6'b000000;
12'b010010011111: data = 6'b010101;
12'b010010100000: data = 6'b111111;
12'b010010100001: data = 6'b111111;
12'b010010100010: data = 6'b111111;
12'b010010100011: data = 6'b111111;
12'b010010100100: data = 6'b111111;
12'b010010100101: data = 6'b111111;
12'b010010100110: data = 6'b111111;
12'b010010100111: data = 6'b111111;
12'b010010101000: data = 6'b111111;
12'b010010101001: data = 6'b111111;
12'b010010101010: data = 6'b111111;
12'b010010101011: data = 6'b111111;
12'b010010101100: data = 6'b111111;
12'b010010101101: data = 6'b111111;
12'b010010101110: data = 6'b111111;
12'b010010101111: data = 6'b111111;
12'b010010110000: data = 6'b111111;
12'b010010110001: data = 6'b111111;
12'b010010110010: data = 6'b111111;
12'b010010110011: data = 6'b111111;
12'b010010110100: data = 6'b111111;
12'b010010110101: data = 6'b111111;
12'b010010110110: data = 6'b111111;
12'b010010110111: data = 6'b111111;
12'b010010111000: data = 6'b111111;
12'b010010111001: data = 6'b111111;
12'b010010111010: data = 6'b111111;
12'b010010111011: data = 6'b111111;
12'b010010111100: data = 6'b111111;
12'b010010111101: data = 6'b111111;
12'b010010111110: data = 6'b111111;
12'b010010111111: data = 6'b111111;
12'b0100101000000: data = 6'b111111;
12'b0100101000001: data = 6'b111111;
12'b0100101000010: data = 6'b111111;
12'b0100101000011: data = 6'b111111;
12'b0100101000100: data = 6'b111111;
12'b0100101000101: data = 6'b111111;
12'b0100101000110: data = 6'b111111;
12'b0100101000111: data = 6'b111111;
12'b0100101001000: data = 6'b111111;
12'b0100101001001: data = 6'b111111;
12'b0100101001010: data = 6'b111111;
12'b0100101001011: data = 6'b111111;
12'b0100101001100: data = 6'b111111;
12'b0100101001101: data = 6'b111111;
12'b0100101001110: data = 6'b111111;
12'b0100101001111: data = 6'b111111;
12'b0100101010000: data = 6'b111111;
12'b0100101010001: data = 6'b111111;
12'b0100101010010: data = 6'b111111;
12'b0100101010011: data = 6'b111111;
12'b0100101010100: data = 6'b111111;
12'b0100101010101: data = 6'b111111;
12'b0100101010110: data = 6'b111111;
12'b0100101010111: data = 6'b111111;
12'b0100101011000: data = 6'b111111;
12'b0100101011001: data = 6'b111111;
12'b0100101011010: data = 6'b111111;
12'b0100101011011: data = 6'b111111;
12'b0100101011100: data = 6'b111111;
12'b0100101011101: data = 6'b111111;
12'b0100101011110: data = 6'b111111;
12'b0100101011111: data = 6'b111111;
12'b0100101100000: data = 6'b111111;
12'b0100101100001: data = 6'b111111;
12'b0100101100010: data = 6'b111111;
12'b0100101100011: data = 6'b111111;
12'b0100101100100: data = 6'b111111;
12'b0100101100101: data = 6'b111111;
12'b0100101100110: data = 6'b111111;
12'b0100101100111: data = 6'b111111;
12'b0100101101000: data = 6'b111111;
12'b0100101101001: data = 6'b111111;
12'b0100101101010: data = 6'b111111;
12'b0100101101011: data = 6'b111111;
12'b0100101101100: data = 6'b111111;
12'b0100101101101: data = 6'b111111;
12'b0100101101110: data = 6'b111111;
12'b0100101101111: data = 6'b111111;
12'b0100101110000: data = 6'b111111;
12'b0100101110001: data = 6'b111111;
12'b0100101110010: data = 6'b111111;
12'b0100101110011: data = 6'b111111;
12'b0100101110100: data = 6'b111111;
12'b0100101110101: data = 6'b111111;
12'b0100101110110: data = 6'b111111;
12'b0100101110111: data = 6'b111111;
12'b0100101111000: data = 6'b111111;
12'b0100101111001: data = 6'b111111;
12'b0100101111010: data = 6'b111111;
12'b0100101111011: data = 6'b111111;
12'b0100101111100: data = 6'b111111;
12'b0100101111101: data = 6'b111111;
12'b0100101111110: data = 6'b111111;
12'b0100101111111: data = 6'b111111;
12'b01001010000000: data = 6'b111111;
12'b01001010000001: data = 6'b111111;
12'b01001010000010: data = 6'b111111;
12'b01001010000011: data = 6'b111111;
12'b01001010000100: data = 6'b111111;
12'b01001010000101: data = 6'b111111;
12'b01001010000110: data = 6'b111111;
12'b01001010000111: data = 6'b111111;
12'b01001010001000: data = 6'b111111;
12'b01001010001001: data = 6'b111111;
12'b01001010001010: data = 6'b111111;
12'b01001010001011: data = 6'b010101;
12'b01001010001100: data = 6'b000000;
12'b01001010001101: data = 6'b000000;
12'b01001010001110: data = 6'b101001;
12'b01001010001111: data = 6'b101010;
12'b01001010010000: data = 6'b101010;
12'b01001010010001: data = 6'b101010;
12'b01001010010010: data = 6'b010101;
12'b01001010010011: data = 6'b010101;
12'b01001010010100: data = 6'b010101;
12'b01001010010101: data = 6'b010101;
12'b01001010010110: data = 6'b010101;
12'b01001010010111: data = 6'b010101;
12'b01001010011000: data = 6'b010101;
12'b01001010011001: data = 6'b010101;
12'b01001010011010: data = 6'b010101;
12'b01001010011011: data = 6'b010101;
12'b01001010011100: data = 6'b010101;
12'b01001010011101: data = 6'b010101;
12'b01001010011110: data = 6'b010101;
12'b01001010011111: data = 6'b010101;
12'b01001010100000: data = 6'b010101;
12'b01001010100001: data = 6'b010101;
12'b01001010100010: data = 6'b010101;
12'b01001010100011: data = 6'b010101;
12'b01001010100100: data = 6'b010101;
12'b01001010100101: data = 6'b010101;
12'b01001010100110: data = 6'b010101;
12'b01001010100111: data = 6'b010101;
12'b01001010101000: data = 6'b010101;
12'b01001010101001: data = 6'b010101;
12'b01001010101010: data = 6'b010101;
12'b010011000000: data = 6'b010101;
12'b010011000001: data = 6'b010101;
12'b010011000010: data = 6'b010101;
12'b010011000011: data = 6'b010101;
12'b010011000100: data = 6'b010101;
12'b010011000101: data = 6'b010101;
12'b010011000110: data = 6'b010101;
12'b010011000111: data = 6'b010101;
12'b010011001000: data = 6'b010101;
12'b010011001001: data = 6'b010101;
12'b010011001010: data = 6'b010101;
12'b010011001011: data = 6'b010101;
12'b010011001100: data = 6'b010101;
12'b010011001101: data = 6'b010101;
12'b010011001110: data = 6'b010101;
12'b010011001111: data = 6'b010101;
12'b010011010000: data = 6'b010101;
12'b010011010001: data = 6'b010101;
12'b010011010010: data = 6'b010101;
12'b010011010011: data = 6'b010101;
12'b010011010100: data = 6'b010101;
12'b010011010101: data = 6'b010101;
12'b010011010110: data = 6'b010101;
12'b010011010111: data = 6'b010101;
12'b010011011000: data = 6'b010101;
12'b010011011001: data = 6'b101010;
12'b010011011010: data = 6'b101010;
12'b010011011011: data = 6'b101010;
12'b010011011100: data = 6'b010101;
12'b010011011101: data = 6'b000000;
12'b010011011110: data = 6'b000000;
12'b010011011111: data = 6'b010101;
12'b010011100000: data = 6'b111111;
12'b010011100001: data = 6'b111111;
12'b010011100010: data = 6'b111111;
12'b010011100011: data = 6'b111111;
12'b010011100100: data = 6'b111111;
12'b010011100101: data = 6'b111111;
12'b010011100110: data = 6'b111111;
12'b010011100111: data = 6'b111111;
12'b010011101000: data = 6'b111111;
12'b010011101001: data = 6'b111111;
12'b010011101010: data = 6'b111111;
12'b010011101011: data = 6'b111111;
12'b010011101100: data = 6'b111111;
12'b010011101101: data = 6'b111111;
12'b010011101110: data = 6'b111111;
12'b010011101111: data = 6'b111111;
12'b010011110000: data = 6'b111111;
12'b010011110001: data = 6'b111111;
12'b010011110010: data = 6'b111111;
12'b010011110011: data = 6'b111111;
12'b010011110100: data = 6'b111111;
12'b010011110101: data = 6'b111111;
12'b010011110110: data = 6'b111111;
12'b010011110111: data = 6'b111111;
12'b010011111000: data = 6'b111111;
12'b010011111001: data = 6'b111111;
12'b010011111010: data = 6'b111111;
12'b010011111011: data = 6'b111111;
12'b010011111100: data = 6'b111111;
12'b010011111101: data = 6'b111111;
12'b010011111110: data = 6'b111111;
12'b010011111111: data = 6'b111111;
12'b0100111000000: data = 6'b111111;
12'b0100111000001: data = 6'b111111;
12'b0100111000010: data = 6'b111111;
12'b0100111000011: data = 6'b111111;
12'b0100111000100: data = 6'b111111;
12'b0100111000101: data = 6'b111111;
12'b0100111000110: data = 6'b111111;
12'b0100111000111: data = 6'b111111;
12'b0100111001000: data = 6'b111111;
12'b0100111001001: data = 6'b111111;
12'b0100111001010: data = 6'b111111;
12'b0100111001011: data = 6'b111111;
12'b0100111001100: data = 6'b111111;
12'b0100111001101: data = 6'b111111;
12'b0100111001110: data = 6'b111111;
12'b0100111001111: data = 6'b111111;
12'b0100111010000: data = 6'b111111;
12'b0100111010001: data = 6'b111111;
12'b0100111010010: data = 6'b111111;
12'b0100111010011: data = 6'b111111;
12'b0100111010100: data = 6'b111111;
12'b0100111010101: data = 6'b111111;
12'b0100111010110: data = 6'b111111;
12'b0100111010111: data = 6'b111111;
12'b0100111011000: data = 6'b111111;
12'b0100111011001: data = 6'b111111;
12'b0100111011010: data = 6'b111111;
12'b0100111011011: data = 6'b111111;
12'b0100111011100: data = 6'b111111;
12'b0100111011101: data = 6'b111111;
12'b0100111011110: data = 6'b111111;
12'b0100111011111: data = 6'b111111;
12'b0100111100000: data = 6'b111111;
12'b0100111100001: data = 6'b111111;
12'b0100111100010: data = 6'b111111;
12'b0100111100011: data = 6'b111111;
12'b0100111100100: data = 6'b111111;
12'b0100111100101: data = 6'b111111;
12'b0100111100110: data = 6'b111111;
12'b0100111100111: data = 6'b111111;
12'b0100111101000: data = 6'b111111;
12'b0100111101001: data = 6'b111111;
12'b0100111101010: data = 6'b111111;
12'b0100111101011: data = 6'b111111;
12'b0100111101100: data = 6'b111111;
12'b0100111101101: data = 6'b111111;
12'b0100111101110: data = 6'b111111;
12'b0100111101111: data = 6'b111111;
12'b0100111110000: data = 6'b111111;
12'b0100111110001: data = 6'b111111;
12'b0100111110010: data = 6'b111111;
12'b0100111110011: data = 6'b111111;
12'b0100111110100: data = 6'b111111;
12'b0100111110101: data = 6'b111111;
12'b0100111110110: data = 6'b111111;
12'b0100111110111: data = 6'b111111;
12'b0100111111000: data = 6'b111111;
12'b0100111111001: data = 6'b111111;
12'b0100111111010: data = 6'b111111;
12'b0100111111011: data = 6'b111111;
12'b0100111111100: data = 6'b111111;
12'b0100111111101: data = 6'b111111;
12'b0100111111110: data = 6'b111111;
12'b0100111111111: data = 6'b111111;
12'b01001110000000: data = 6'b111111;
12'b01001110000001: data = 6'b111111;
12'b01001110000010: data = 6'b111111;
12'b01001110000011: data = 6'b111111;
12'b01001110000100: data = 6'b111111;
12'b01001110000101: data = 6'b111111;
12'b01001110000110: data = 6'b111111;
12'b01001110000111: data = 6'b111111;
12'b01001110001000: data = 6'b111111;
12'b01001110001001: data = 6'b111111;
12'b01001110001010: data = 6'b111111;
12'b01001110001011: data = 6'b010101;
12'b01001110001100: data = 6'b000000;
12'b01001110001101: data = 6'b000000;
12'b01001110001110: data = 6'b101001;
12'b01001110001111: data = 6'b101010;
12'b01001110010000: data = 6'b101010;
12'b01001110010001: data = 6'b101010;
12'b01001110010010: data = 6'b010101;
12'b01001110010011: data = 6'b010101;
12'b01001110010100: data = 6'b010101;
12'b01001110010101: data = 6'b010101;
12'b01001110010110: data = 6'b010101;
12'b01001110010111: data = 6'b010101;
12'b01001110011000: data = 6'b010101;
12'b01001110011001: data = 6'b010101;
12'b01001110011010: data = 6'b010101;
12'b01001110011011: data = 6'b010101;
12'b01001110011100: data = 6'b010101;
12'b01001110011101: data = 6'b010101;
12'b01001110011110: data = 6'b010101;
12'b01001110011111: data = 6'b010101;
12'b01001110100000: data = 6'b010101;
12'b01001110100001: data = 6'b010101;
12'b01001110100010: data = 6'b010101;
12'b01001110100011: data = 6'b010101;
12'b01001110100100: data = 6'b010101;
12'b01001110100101: data = 6'b010101;
12'b01001110100110: data = 6'b010101;
12'b01001110100111: data = 6'b010101;
12'b01001110101000: data = 6'b010101;
12'b01001110101001: data = 6'b010101;
12'b01001110101010: data = 6'b010101;
12'b010100000000: data = 6'b010101;
12'b010100000001: data = 6'b010101;
12'b010100000010: data = 6'b010101;
12'b010100000011: data = 6'b010101;
12'b010100000100: data = 6'b010101;
12'b010100000101: data = 6'b010101;
12'b010100000110: data = 6'b010101;
12'b010100000111: data = 6'b010101;
12'b010100001000: data = 6'b010101;
12'b010100001001: data = 6'b010101;
12'b010100001010: data = 6'b010101;
12'b010100001011: data = 6'b010101;
12'b010100001100: data = 6'b010101;
12'b010100001101: data = 6'b010101;
12'b010100001110: data = 6'b010101;
12'b010100001111: data = 6'b010101;
12'b010100010000: data = 6'b010101;
12'b010100010001: data = 6'b010101;
12'b010100010010: data = 6'b010101;
12'b010100010011: data = 6'b010101;
12'b010100010100: data = 6'b010101;
12'b010100010101: data = 6'b010101;
12'b010100010110: data = 6'b010101;
12'b010100010111: data = 6'b010101;
12'b010100011000: data = 6'b010101;
12'b010100011001: data = 6'b101010;
12'b010100011010: data = 6'b101010;
12'b010100011011: data = 6'b101010;
12'b010100011100: data = 6'b010101;
12'b010100011101: data = 6'b000000;
12'b010100011110: data = 6'b000000;
12'b010100011111: data = 6'b010101;
12'b010100100000: data = 6'b111111;
12'b010100100001: data = 6'b111111;
12'b010100100010: data = 6'b111111;
12'b010100100011: data = 6'b111111;
12'b010100100100: data = 6'b111111;
12'b010100100101: data = 6'b111111;
12'b010100100110: data = 6'b111111;
12'b010100100111: data = 6'b111111;
12'b010100101000: data = 6'b111111;
12'b010100101001: data = 6'b111111;
12'b010100101010: data = 6'b111111;
12'b010100101011: data = 6'b111111;
12'b010100101100: data = 6'b111111;
12'b010100101101: data = 6'b111111;
12'b010100101110: data = 6'b111111;
12'b010100101111: data = 6'b111111;
12'b010100110000: data = 6'b111111;
12'b010100110001: data = 6'b111111;
12'b010100110010: data = 6'b111111;
12'b010100110011: data = 6'b111111;
12'b010100110100: data = 6'b111111;
12'b010100110101: data = 6'b111111;
12'b010100110110: data = 6'b111111;
12'b010100110111: data = 6'b111111;
12'b010100111000: data = 6'b111111;
12'b010100111001: data = 6'b111111;
12'b010100111010: data = 6'b111111;
12'b010100111011: data = 6'b111111;
12'b010100111100: data = 6'b111111;
12'b010100111101: data = 6'b111111;
12'b010100111110: data = 6'b111111;
12'b010100111111: data = 6'b111111;
12'b0101001000000: data = 6'b111111;
12'b0101001000001: data = 6'b111111;
12'b0101001000010: data = 6'b111111;
12'b0101001000011: data = 6'b111111;
12'b0101001000100: data = 6'b111111;
12'b0101001000101: data = 6'b111111;
12'b0101001000110: data = 6'b111111;
12'b0101001000111: data = 6'b111111;
12'b0101001001000: data = 6'b111111;
12'b0101001001001: data = 6'b111111;
12'b0101001001010: data = 6'b111111;
12'b0101001001011: data = 6'b111111;
12'b0101001001100: data = 6'b111111;
12'b0101001001101: data = 6'b111111;
12'b0101001001110: data = 6'b111111;
12'b0101001001111: data = 6'b111111;
12'b0101001010000: data = 6'b111111;
12'b0101001010001: data = 6'b111111;
12'b0101001010010: data = 6'b111111;
12'b0101001010011: data = 6'b111111;
12'b0101001010100: data = 6'b111111;
12'b0101001010101: data = 6'b111111;
12'b0101001010110: data = 6'b111111;
12'b0101001010111: data = 6'b111111;
12'b0101001011000: data = 6'b111111;
12'b0101001011001: data = 6'b111111;
12'b0101001011010: data = 6'b111111;
12'b0101001011011: data = 6'b111111;
12'b0101001011100: data = 6'b111111;
12'b0101001011101: data = 6'b111111;
12'b0101001011110: data = 6'b111111;
12'b0101001011111: data = 6'b111111;
12'b0101001100000: data = 6'b111111;
12'b0101001100001: data = 6'b111111;
12'b0101001100010: data = 6'b111111;
12'b0101001100011: data = 6'b111111;
12'b0101001100100: data = 6'b111111;
12'b0101001100101: data = 6'b111111;
12'b0101001100110: data = 6'b111111;
12'b0101001100111: data = 6'b111111;
12'b0101001101000: data = 6'b111111;
12'b0101001101001: data = 6'b111111;
12'b0101001101010: data = 6'b111111;
12'b0101001101011: data = 6'b111111;
12'b0101001101100: data = 6'b111111;
12'b0101001101101: data = 6'b111111;
12'b0101001101110: data = 6'b111111;
12'b0101001101111: data = 6'b111111;
12'b0101001110000: data = 6'b111111;
12'b0101001110001: data = 6'b111111;
12'b0101001110010: data = 6'b111111;
12'b0101001110011: data = 6'b111111;
12'b0101001110100: data = 6'b111111;
12'b0101001110101: data = 6'b111111;
12'b0101001110110: data = 6'b111111;
12'b0101001110111: data = 6'b111111;
12'b0101001111000: data = 6'b111111;
12'b0101001111001: data = 6'b111111;
12'b0101001111010: data = 6'b111111;
12'b0101001111011: data = 6'b111111;
12'b0101001111100: data = 6'b111111;
12'b0101001111101: data = 6'b111111;
12'b0101001111110: data = 6'b111111;
12'b0101001111111: data = 6'b111111;
12'b01010010000000: data = 6'b111111;
12'b01010010000001: data = 6'b111111;
12'b01010010000010: data = 6'b111111;
12'b01010010000011: data = 6'b111111;
12'b01010010000100: data = 6'b111111;
12'b01010010000101: data = 6'b111111;
12'b01010010000110: data = 6'b111111;
12'b01010010000111: data = 6'b111111;
12'b01010010001000: data = 6'b111111;
12'b01010010001001: data = 6'b111111;
12'b01010010001010: data = 6'b111111;
12'b01010010001011: data = 6'b010101;
12'b01010010001100: data = 6'b000000;
12'b01010010001101: data = 6'b000000;
12'b01010010001110: data = 6'b101001;
12'b01010010001111: data = 6'b101010;
12'b01010010010000: data = 6'b101010;
12'b01010010010001: data = 6'b101010;
12'b01010010010010: data = 6'b010101;
12'b01010010010011: data = 6'b010101;
12'b01010010010100: data = 6'b010101;
12'b01010010010101: data = 6'b010101;
12'b01010010010110: data = 6'b010101;
12'b01010010010111: data = 6'b010101;
12'b01010010011000: data = 6'b010101;
12'b01010010011001: data = 6'b010101;
12'b01010010011010: data = 6'b010101;
12'b01010010011011: data = 6'b010101;
12'b01010010011100: data = 6'b010101;
12'b01010010011101: data = 6'b010101;
12'b01010010011110: data = 6'b010101;
12'b01010010011111: data = 6'b010101;
12'b01010010100000: data = 6'b010101;
12'b01010010100001: data = 6'b010101;
12'b01010010100010: data = 6'b010101;
12'b01010010100011: data = 6'b010101;
12'b01010010100100: data = 6'b010101;
12'b01010010100101: data = 6'b010101;
12'b01010010100110: data = 6'b010101;
12'b01010010100111: data = 6'b010101;
12'b01010010101000: data = 6'b010101;
12'b01010010101001: data = 6'b010101;
12'b01010010101010: data = 6'b010101;
12'b010101000000: data = 6'b010101;
12'b010101000001: data = 6'b010101;
12'b010101000010: data = 6'b010101;
12'b010101000011: data = 6'b010101;
12'b010101000100: data = 6'b010101;
12'b010101000101: data = 6'b010101;
12'b010101000110: data = 6'b010101;
12'b010101000111: data = 6'b010101;
12'b010101001000: data = 6'b010101;
12'b010101001001: data = 6'b010101;
12'b010101001010: data = 6'b010101;
12'b010101001011: data = 6'b010101;
12'b010101001100: data = 6'b010101;
12'b010101001101: data = 6'b010101;
12'b010101001110: data = 6'b010101;
12'b010101001111: data = 6'b010101;
12'b010101010000: data = 6'b010101;
12'b010101010001: data = 6'b010101;
12'b010101010010: data = 6'b010101;
12'b010101010011: data = 6'b010101;
12'b010101010100: data = 6'b010101;
12'b010101010101: data = 6'b010101;
12'b010101010110: data = 6'b010101;
12'b010101010111: data = 6'b010101;
12'b010101011000: data = 6'b010101;
12'b010101011001: data = 6'b101010;
12'b010101011010: data = 6'b101010;
12'b010101011011: data = 6'b101010;
12'b010101011100: data = 6'b010101;
12'b010101011101: data = 6'b000000;
12'b010101011110: data = 6'b000000;
12'b010101011111: data = 6'b010101;
12'b010101100000: data = 6'b111111;
12'b010101100001: data = 6'b111111;
12'b010101100010: data = 6'b111111;
12'b010101100011: data = 6'b111111;
12'b010101100100: data = 6'b111111;
12'b010101100101: data = 6'b111111;
12'b010101100110: data = 6'b111111;
12'b010101100111: data = 6'b111111;
12'b010101101000: data = 6'b111111;
12'b010101101001: data = 6'b111111;
12'b010101101010: data = 6'b111111;
12'b010101101011: data = 6'b111111;
12'b010101101100: data = 6'b111111;
12'b010101101101: data = 6'b111111;
12'b010101101110: data = 6'b111111;
12'b010101101111: data = 6'b111111;
12'b010101110000: data = 6'b111111;
12'b010101110001: data = 6'b111111;
12'b010101110010: data = 6'b111111;
12'b010101110011: data = 6'b111111;
12'b010101110100: data = 6'b111111;
12'b010101110101: data = 6'b111111;
12'b010101110110: data = 6'b111111;
12'b010101110111: data = 6'b111111;
12'b010101111000: data = 6'b111111;
12'b010101111001: data = 6'b111111;
12'b010101111010: data = 6'b111111;
12'b010101111011: data = 6'b111111;
12'b010101111100: data = 6'b111111;
12'b010101111101: data = 6'b111111;
12'b010101111110: data = 6'b111111;
12'b010101111111: data = 6'b111111;
12'b0101011000000: data = 6'b111111;
12'b0101011000001: data = 6'b111111;
12'b0101011000010: data = 6'b111111;
12'b0101011000011: data = 6'b111111;
12'b0101011000100: data = 6'b111111;
12'b0101011000101: data = 6'b111111;
12'b0101011000110: data = 6'b111111;
12'b0101011000111: data = 6'b111111;
12'b0101011001000: data = 6'b111111;
12'b0101011001001: data = 6'b111111;
12'b0101011001010: data = 6'b111111;
12'b0101011001011: data = 6'b111111;
12'b0101011001100: data = 6'b111111;
12'b0101011001101: data = 6'b111111;
12'b0101011001110: data = 6'b111111;
12'b0101011001111: data = 6'b111111;
12'b0101011010000: data = 6'b111111;
12'b0101011010001: data = 6'b111111;
12'b0101011010010: data = 6'b111111;
12'b0101011010011: data = 6'b111111;
12'b0101011010100: data = 6'b111111;
12'b0101011010101: data = 6'b111111;
12'b0101011010110: data = 6'b111111;
12'b0101011010111: data = 6'b111111;
12'b0101011011000: data = 6'b111111;
12'b0101011011001: data = 6'b111111;
12'b0101011011010: data = 6'b111111;
12'b0101011011011: data = 6'b111111;
12'b0101011011100: data = 6'b111111;
12'b0101011011101: data = 6'b111111;
12'b0101011011110: data = 6'b111111;
12'b0101011011111: data = 6'b111111;
12'b0101011100000: data = 6'b111111;
12'b0101011100001: data = 6'b111111;
12'b0101011100010: data = 6'b111111;
12'b0101011100011: data = 6'b111111;
12'b0101011100100: data = 6'b111111;
12'b0101011100101: data = 6'b111111;
12'b0101011100110: data = 6'b111111;
12'b0101011100111: data = 6'b111111;
12'b0101011101000: data = 6'b111111;
12'b0101011101001: data = 6'b111111;
12'b0101011101010: data = 6'b111111;
12'b0101011101011: data = 6'b111111;
12'b0101011101100: data = 6'b111111;
12'b0101011101101: data = 6'b111111;
12'b0101011101110: data = 6'b111111;
12'b0101011101111: data = 6'b111111;
12'b0101011110000: data = 6'b111111;
12'b0101011110001: data = 6'b111111;
12'b0101011110010: data = 6'b111111;
12'b0101011110011: data = 6'b111111;
12'b0101011110100: data = 6'b111111;
12'b0101011110101: data = 6'b111111;
12'b0101011110110: data = 6'b111111;
12'b0101011110111: data = 6'b111111;
12'b0101011111000: data = 6'b111111;
12'b0101011111001: data = 6'b111111;
12'b0101011111010: data = 6'b111111;
12'b0101011111011: data = 6'b111111;
12'b0101011111100: data = 6'b111111;
12'b0101011111101: data = 6'b111111;
12'b0101011111110: data = 6'b111111;
12'b0101011111111: data = 6'b111111;
12'b01010110000000: data = 6'b111111;
12'b01010110000001: data = 6'b111111;
12'b01010110000010: data = 6'b111111;
12'b01010110000011: data = 6'b111111;
12'b01010110000100: data = 6'b111111;
12'b01010110000101: data = 6'b111111;
12'b01010110000110: data = 6'b111111;
12'b01010110000111: data = 6'b111111;
12'b01010110001000: data = 6'b111111;
12'b01010110001001: data = 6'b111111;
12'b01010110001010: data = 6'b111111;
12'b01010110001011: data = 6'b010101;
12'b01010110001100: data = 6'b000000;
12'b01010110001101: data = 6'b000000;
12'b01010110001110: data = 6'b101001;
12'b01010110001111: data = 6'b101010;
12'b01010110010000: data = 6'b101010;
12'b01010110010001: data = 6'b101010;
12'b01010110010010: data = 6'b010101;
12'b01010110010011: data = 6'b010101;
12'b01010110010100: data = 6'b010101;
12'b01010110010101: data = 6'b010101;
12'b01010110010110: data = 6'b010101;
12'b01010110010111: data = 6'b010101;
12'b01010110011000: data = 6'b010101;
12'b01010110011001: data = 6'b010101;
12'b01010110011010: data = 6'b010101;
12'b01010110011011: data = 6'b010101;
12'b01010110011100: data = 6'b010101;
12'b01010110011101: data = 6'b010101;
12'b01010110011110: data = 6'b010101;
12'b01010110011111: data = 6'b010101;
12'b01010110100000: data = 6'b010101;
12'b01010110100001: data = 6'b010101;
12'b01010110100010: data = 6'b010101;
12'b01010110100011: data = 6'b010101;
12'b01010110100100: data = 6'b010101;
12'b01010110100101: data = 6'b010101;
12'b01010110100110: data = 6'b010101;
12'b01010110100111: data = 6'b010101;
12'b01010110101000: data = 6'b010101;
12'b01010110101001: data = 6'b010101;
12'b01010110101010: data = 6'b010101;
12'b010110000000: data = 6'b010101;
12'b010110000001: data = 6'b010101;
12'b010110000010: data = 6'b010101;
12'b010110000011: data = 6'b010101;
12'b010110000100: data = 6'b010101;
12'b010110000101: data = 6'b010101;
12'b010110000110: data = 6'b010101;
12'b010110000111: data = 6'b010101;
12'b010110001000: data = 6'b010101;
12'b010110001001: data = 6'b010101;
12'b010110001010: data = 6'b010101;
12'b010110001011: data = 6'b010101;
12'b010110001100: data = 6'b010101;
12'b010110001101: data = 6'b010101;
12'b010110001110: data = 6'b010101;
12'b010110001111: data = 6'b010101;
12'b010110010000: data = 6'b010101;
12'b010110010001: data = 6'b010101;
12'b010110010010: data = 6'b010101;
12'b010110010011: data = 6'b010101;
12'b010110010100: data = 6'b010101;
12'b010110010101: data = 6'b010101;
12'b010110010110: data = 6'b010101;
12'b010110010111: data = 6'b010101;
12'b010110011000: data = 6'b010101;
12'b010110011001: data = 6'b101010;
12'b010110011010: data = 6'b101010;
12'b010110011011: data = 6'b101010;
12'b010110011100: data = 6'b010101;
12'b010110011101: data = 6'b000000;
12'b010110011110: data = 6'b000000;
12'b010110011111: data = 6'b010101;
12'b010110100000: data = 6'b111111;
12'b010110100001: data = 6'b111111;
12'b010110100010: data = 6'b111111;
12'b010110100011: data = 6'b111111;
12'b010110100100: data = 6'b111111;
12'b010110100101: data = 6'b111111;
12'b010110100110: data = 6'b111111;
12'b010110100111: data = 6'b111111;
12'b010110101000: data = 6'b111111;
12'b010110101001: data = 6'b111111;
12'b010110101010: data = 6'b111111;
12'b010110101011: data = 6'b111111;
12'b010110101100: data = 6'b111111;
12'b010110101101: data = 6'b111111;
12'b010110101110: data = 6'b111111;
12'b010110101111: data = 6'b111111;
12'b010110110000: data = 6'b111111;
12'b010110110001: data = 6'b111111;
12'b010110110010: data = 6'b111111;
12'b010110110011: data = 6'b111111;
12'b010110110100: data = 6'b111111;
12'b010110110101: data = 6'b111111;
12'b010110110110: data = 6'b111111;
12'b010110110111: data = 6'b111111;
12'b010110111000: data = 6'b111111;
12'b010110111001: data = 6'b111111;
12'b010110111010: data = 6'b111111;
12'b010110111011: data = 6'b111111;
12'b010110111100: data = 6'b111111;
12'b010110111101: data = 6'b111111;
12'b010110111110: data = 6'b111111;
12'b010110111111: data = 6'b111111;
12'b0101101000000: data = 6'b111111;
12'b0101101000001: data = 6'b111111;
12'b0101101000010: data = 6'b111111;
12'b0101101000011: data = 6'b111111;
12'b0101101000100: data = 6'b111111;
12'b0101101000101: data = 6'b111111;
12'b0101101000110: data = 6'b111111;
12'b0101101000111: data = 6'b111111;
12'b0101101001000: data = 6'b111111;
12'b0101101001001: data = 6'b111111;
12'b0101101001010: data = 6'b111111;
12'b0101101001011: data = 6'b111111;
12'b0101101001100: data = 6'b111111;
12'b0101101001101: data = 6'b111111;
12'b0101101001110: data = 6'b111111;
12'b0101101001111: data = 6'b111111;
12'b0101101010000: data = 6'b111111;
12'b0101101010001: data = 6'b111111;
12'b0101101010010: data = 6'b111111;
12'b0101101010011: data = 6'b111111;
12'b0101101010100: data = 6'b111111;
12'b0101101010101: data = 6'b111111;
12'b0101101010110: data = 6'b111111;
12'b0101101010111: data = 6'b111111;
12'b0101101011000: data = 6'b111111;
12'b0101101011001: data = 6'b111111;
12'b0101101011010: data = 6'b111111;
12'b0101101011011: data = 6'b111111;
12'b0101101011100: data = 6'b111111;
12'b0101101011101: data = 6'b111111;
12'b0101101011110: data = 6'b111111;
12'b0101101011111: data = 6'b111111;
12'b0101101100000: data = 6'b111111;
12'b0101101100001: data = 6'b111111;
12'b0101101100010: data = 6'b111111;
12'b0101101100011: data = 6'b111111;
12'b0101101100100: data = 6'b111111;
12'b0101101100101: data = 6'b111111;
12'b0101101100110: data = 6'b111111;
12'b0101101100111: data = 6'b111111;
12'b0101101101000: data = 6'b111111;
12'b0101101101001: data = 6'b111111;
12'b0101101101010: data = 6'b111111;
12'b0101101101011: data = 6'b111111;
12'b0101101101100: data = 6'b111111;
12'b0101101101101: data = 6'b111111;
12'b0101101101110: data = 6'b111111;
12'b0101101101111: data = 6'b111111;
12'b0101101110000: data = 6'b111111;
12'b0101101110001: data = 6'b111111;
12'b0101101110010: data = 6'b111111;
12'b0101101110011: data = 6'b111111;
12'b0101101110100: data = 6'b111111;
12'b0101101110101: data = 6'b111111;
12'b0101101110110: data = 6'b111111;
12'b0101101110111: data = 6'b111111;
12'b0101101111000: data = 6'b111111;
12'b0101101111001: data = 6'b111111;
12'b0101101111010: data = 6'b111111;
12'b0101101111011: data = 6'b111111;
12'b0101101111100: data = 6'b111111;
12'b0101101111101: data = 6'b111111;
12'b0101101111110: data = 6'b111111;
12'b0101101111111: data = 6'b111111;
12'b01011010000000: data = 6'b111111;
12'b01011010000001: data = 6'b111111;
12'b01011010000010: data = 6'b111111;
12'b01011010000011: data = 6'b111111;
12'b01011010000100: data = 6'b111111;
12'b01011010000101: data = 6'b111111;
12'b01011010000110: data = 6'b111111;
12'b01011010000111: data = 6'b111111;
12'b01011010001000: data = 6'b111111;
12'b01011010001001: data = 6'b111111;
12'b01011010001010: data = 6'b111111;
12'b01011010001011: data = 6'b010101;
12'b01011010001100: data = 6'b000000;
12'b01011010001101: data = 6'b000000;
12'b01011010001110: data = 6'b101010;
12'b01011010001111: data = 6'b101010;
12'b01011010010000: data = 6'b101010;
12'b01011010010001: data = 6'b101010;
12'b01011010010010: data = 6'b010101;
12'b01011010010011: data = 6'b010101;
12'b01011010010100: data = 6'b010101;
12'b01011010010101: data = 6'b010101;
12'b01011010010110: data = 6'b010101;
12'b01011010010111: data = 6'b010101;
12'b01011010011000: data = 6'b010101;
12'b01011010011001: data = 6'b010101;
12'b01011010011010: data = 6'b010101;
12'b01011010011011: data = 6'b010101;
12'b01011010011100: data = 6'b010101;
12'b01011010011101: data = 6'b010101;
12'b01011010011110: data = 6'b010101;
12'b01011010011111: data = 6'b010101;
12'b01011010100000: data = 6'b010101;
12'b01011010100001: data = 6'b010101;
12'b01011010100010: data = 6'b010101;
12'b01011010100011: data = 6'b010101;
12'b01011010100100: data = 6'b010101;
12'b01011010100101: data = 6'b010101;
12'b01011010100110: data = 6'b010101;
12'b01011010100111: data = 6'b010101;
12'b01011010101000: data = 6'b010101;
12'b01011010101001: data = 6'b010101;
12'b01011010101010: data = 6'b010101;
12'b010111000000: data = 6'b010101;
12'b010111000001: data = 6'b010101;
12'b010111000010: data = 6'b010101;
12'b010111000011: data = 6'b010101;
12'b010111000100: data = 6'b010101;
12'b010111000101: data = 6'b010101;
12'b010111000110: data = 6'b010101;
12'b010111000111: data = 6'b010101;
12'b010111001000: data = 6'b010101;
12'b010111001001: data = 6'b010101;
12'b010111001010: data = 6'b010101;
12'b010111001011: data = 6'b010101;
12'b010111001100: data = 6'b010101;
12'b010111001101: data = 6'b010101;
12'b010111001110: data = 6'b010101;
12'b010111001111: data = 6'b010101;
12'b010111010000: data = 6'b010101;
12'b010111010001: data = 6'b010101;
12'b010111010010: data = 6'b010101;
12'b010111010011: data = 6'b010101;
12'b010111010100: data = 6'b010101;
12'b010111010101: data = 6'b010101;
12'b010111010110: data = 6'b010101;
12'b010111010111: data = 6'b010101;
12'b010111011000: data = 6'b010101;
12'b010111011001: data = 6'b101010;
12'b010111011010: data = 6'b101010;
12'b010111011011: data = 6'b101010;
12'b010111011100: data = 6'b010101;
12'b010111011101: data = 6'b000000;
12'b010111011110: data = 6'b000000;
12'b010111011111: data = 6'b010101;
12'b010111100000: data = 6'b111111;
12'b010111100001: data = 6'b111111;
12'b010111100010: data = 6'b111111;
12'b010111100011: data = 6'b111111;
12'b010111100100: data = 6'b111111;
12'b010111100101: data = 6'b111111;
12'b010111100110: data = 6'b111111;
12'b010111100111: data = 6'b111111;
12'b010111101000: data = 6'b111111;
12'b010111101001: data = 6'b111111;
12'b010111101010: data = 6'b111111;
12'b010111101011: data = 6'b111111;
12'b010111101100: data = 6'b111111;
12'b010111101101: data = 6'b111111;
12'b010111101110: data = 6'b111111;
12'b010111101111: data = 6'b111111;
12'b010111110000: data = 6'b111111;
12'b010111110001: data = 6'b111111;
12'b010111110010: data = 6'b111111;
12'b010111110011: data = 6'b111111;
12'b010111110100: data = 6'b111111;
12'b010111110101: data = 6'b111111;
12'b010111110110: data = 6'b111111;
12'b010111110111: data = 6'b111111;
12'b010111111000: data = 6'b111111;
12'b010111111001: data = 6'b111111;
12'b010111111010: data = 6'b111111;
12'b010111111011: data = 6'b111111;
12'b010111111100: data = 6'b111111;
12'b010111111101: data = 6'b111111;
12'b010111111110: data = 6'b111111;
12'b010111111111: data = 6'b111111;
12'b0101111000000: data = 6'b111111;
12'b0101111000001: data = 6'b111111;
12'b0101111000010: data = 6'b111111;
12'b0101111000011: data = 6'b111111;
12'b0101111000100: data = 6'b111111;
12'b0101111000101: data = 6'b111111;
12'b0101111000110: data = 6'b111111;
12'b0101111000111: data = 6'b111111;
12'b0101111001000: data = 6'b111111;
12'b0101111001001: data = 6'b111111;
12'b0101111001010: data = 6'b111111;
12'b0101111001011: data = 6'b111111;
12'b0101111001100: data = 6'b111111;
12'b0101111001101: data = 6'b111111;
12'b0101111001110: data = 6'b111111;
12'b0101111001111: data = 6'b111111;
12'b0101111010000: data = 6'b111111;
12'b0101111010001: data = 6'b111111;
12'b0101111010010: data = 6'b111111;
12'b0101111010011: data = 6'b111111;
12'b0101111010100: data = 6'b111111;
12'b0101111010101: data = 6'b111111;
12'b0101111010110: data = 6'b111111;
12'b0101111010111: data = 6'b111111;
12'b0101111011000: data = 6'b111111;
12'b0101111011001: data = 6'b111111;
12'b0101111011010: data = 6'b111111;
12'b0101111011011: data = 6'b111111;
12'b0101111011100: data = 6'b111111;
12'b0101111011101: data = 6'b111111;
12'b0101111011110: data = 6'b111111;
12'b0101111011111: data = 6'b111111;
12'b0101111100000: data = 6'b111111;
12'b0101111100001: data = 6'b111111;
12'b0101111100010: data = 6'b111111;
12'b0101111100011: data = 6'b111111;
12'b0101111100100: data = 6'b111111;
12'b0101111100101: data = 6'b111111;
12'b0101111100110: data = 6'b111111;
12'b0101111100111: data = 6'b111111;
12'b0101111101000: data = 6'b111111;
12'b0101111101001: data = 6'b111111;
12'b0101111101010: data = 6'b111111;
12'b0101111101011: data = 6'b111111;
12'b0101111101100: data = 6'b111111;
12'b0101111101101: data = 6'b111111;
12'b0101111101110: data = 6'b111111;
12'b0101111101111: data = 6'b111111;
12'b0101111110000: data = 6'b111111;
12'b0101111110001: data = 6'b111111;
12'b0101111110010: data = 6'b111111;
12'b0101111110011: data = 6'b111111;
12'b0101111110100: data = 6'b111111;
12'b0101111110101: data = 6'b111111;
12'b0101111110110: data = 6'b111111;
12'b0101111110111: data = 6'b111111;
12'b0101111111000: data = 6'b111111;
12'b0101111111001: data = 6'b111111;
12'b0101111111010: data = 6'b111111;
12'b0101111111011: data = 6'b111111;
12'b0101111111100: data = 6'b111111;
12'b0101111111101: data = 6'b111111;
12'b0101111111110: data = 6'b111111;
12'b0101111111111: data = 6'b111111;
12'b01011110000000: data = 6'b111111;
12'b01011110000001: data = 6'b111111;
12'b01011110000010: data = 6'b111111;
12'b01011110000011: data = 6'b111111;
12'b01011110000100: data = 6'b111111;
12'b01011110000101: data = 6'b111111;
12'b01011110000110: data = 6'b111111;
12'b01011110000111: data = 6'b111111;
12'b01011110001000: data = 6'b111111;
12'b01011110001001: data = 6'b111111;
12'b01011110001010: data = 6'b111111;
12'b01011110001011: data = 6'b010101;
12'b01011110001100: data = 6'b000000;
12'b01011110001101: data = 6'b000000;
12'b01011110001110: data = 6'b101010;
12'b01011110001111: data = 6'b101010;
12'b01011110010000: data = 6'b101010;
12'b01011110010001: data = 6'b101010;
12'b01011110010010: data = 6'b010101;
12'b01011110010011: data = 6'b010101;
12'b01011110010100: data = 6'b010101;
12'b01011110010101: data = 6'b010101;
12'b01011110010110: data = 6'b010101;
12'b01011110010111: data = 6'b010101;
12'b01011110011000: data = 6'b010101;
12'b01011110011001: data = 6'b010101;
12'b01011110011010: data = 6'b010101;
12'b01011110011011: data = 6'b010101;
12'b01011110011100: data = 6'b010101;
12'b01011110011101: data = 6'b010101;
12'b01011110011110: data = 6'b010101;
12'b01011110011111: data = 6'b010101;
12'b01011110100000: data = 6'b010101;
12'b01011110100001: data = 6'b010101;
12'b01011110100010: data = 6'b010101;
12'b01011110100011: data = 6'b010101;
12'b01011110100100: data = 6'b010101;
12'b01011110100101: data = 6'b010101;
12'b01011110100110: data = 6'b010101;
12'b01011110100111: data = 6'b010101;
12'b01011110101000: data = 6'b010101;
12'b01011110101001: data = 6'b010101;
12'b01011110101010: data = 6'b010101;
12'b011000000000: data = 6'b010101;
12'b011000000001: data = 6'b010101;
12'b011000000010: data = 6'b010101;
12'b011000000011: data = 6'b010101;
12'b011000000100: data = 6'b010101;
12'b011000000101: data = 6'b010101;
12'b011000000110: data = 6'b010101;
12'b011000000111: data = 6'b010101;
12'b011000001000: data = 6'b010101;
12'b011000001001: data = 6'b010101;
12'b011000001010: data = 6'b010101;
12'b011000001011: data = 6'b010101;
12'b011000001100: data = 6'b010101;
12'b011000001101: data = 6'b010101;
12'b011000001110: data = 6'b010101;
12'b011000001111: data = 6'b010101;
12'b011000010000: data = 6'b010101;
12'b011000010001: data = 6'b010101;
12'b011000010010: data = 6'b010101;
12'b011000010011: data = 6'b010101;
12'b011000010100: data = 6'b010101;
12'b011000010101: data = 6'b010101;
12'b011000010110: data = 6'b010101;
12'b011000010111: data = 6'b010101;
12'b011000011000: data = 6'b010101;
12'b011000011001: data = 6'b101010;
12'b011000011010: data = 6'b101010;
12'b011000011011: data = 6'b101010;
12'b011000011100: data = 6'b010101;
12'b011000011101: data = 6'b000000;
12'b011000011110: data = 6'b000000;
12'b011000011111: data = 6'b010101;
12'b011000100000: data = 6'b111111;
12'b011000100001: data = 6'b111111;
12'b011000100010: data = 6'b111111;
12'b011000100011: data = 6'b111111;
12'b011000100100: data = 6'b111111;
12'b011000100101: data = 6'b111111;
12'b011000100110: data = 6'b111111;
12'b011000100111: data = 6'b111111;
12'b011000101000: data = 6'b111111;
12'b011000101001: data = 6'b111111;
12'b011000101010: data = 6'b111111;
12'b011000101011: data = 6'b111111;
12'b011000101100: data = 6'b111111;
12'b011000101101: data = 6'b111111;
12'b011000101110: data = 6'b111111;
12'b011000101111: data = 6'b111111;
12'b011000110000: data = 6'b111111;
12'b011000110001: data = 6'b111111;
12'b011000110010: data = 6'b111111;
12'b011000110011: data = 6'b111111;
12'b011000110100: data = 6'b111111;
12'b011000110101: data = 6'b111111;
12'b011000110110: data = 6'b111111;
12'b011000110111: data = 6'b111111;
12'b011000111000: data = 6'b111111;
12'b011000111001: data = 6'b111111;
12'b011000111010: data = 6'b111111;
12'b011000111011: data = 6'b111111;
12'b011000111100: data = 6'b111111;
12'b011000111101: data = 6'b111111;
12'b011000111110: data = 6'b111111;
12'b011000111111: data = 6'b111111;
12'b0110001000000: data = 6'b111111;
12'b0110001000001: data = 6'b111111;
12'b0110001000010: data = 6'b111111;
12'b0110001000011: data = 6'b111111;
12'b0110001000100: data = 6'b111111;
12'b0110001000101: data = 6'b111111;
12'b0110001000110: data = 6'b111111;
12'b0110001000111: data = 6'b111111;
12'b0110001001000: data = 6'b111111;
12'b0110001001001: data = 6'b111111;
12'b0110001001010: data = 6'b111111;
12'b0110001001011: data = 6'b111111;
12'b0110001001100: data = 6'b111111;
12'b0110001001101: data = 6'b111111;
12'b0110001001110: data = 6'b111111;
12'b0110001001111: data = 6'b111111;
12'b0110001010000: data = 6'b111111;
12'b0110001010001: data = 6'b111111;
12'b0110001010010: data = 6'b111111;
12'b0110001010011: data = 6'b111111;
12'b0110001010100: data = 6'b111111;
12'b0110001010101: data = 6'b111111;
12'b0110001010110: data = 6'b111111;
12'b0110001010111: data = 6'b111111;
12'b0110001011000: data = 6'b111111;
12'b0110001011001: data = 6'b111111;
12'b0110001011010: data = 6'b111111;
12'b0110001011011: data = 6'b111111;
12'b0110001011100: data = 6'b111111;
12'b0110001011101: data = 6'b111111;
12'b0110001011110: data = 6'b111111;
12'b0110001011111: data = 6'b111111;
12'b0110001100000: data = 6'b111111;
12'b0110001100001: data = 6'b111111;
12'b0110001100010: data = 6'b111111;
12'b0110001100011: data = 6'b111111;
12'b0110001100100: data = 6'b111111;
12'b0110001100101: data = 6'b111111;
12'b0110001100110: data = 6'b111111;
12'b0110001100111: data = 6'b111111;
12'b0110001101000: data = 6'b111111;
12'b0110001101001: data = 6'b111111;
12'b0110001101010: data = 6'b111111;
12'b0110001101011: data = 6'b111111;
12'b0110001101100: data = 6'b111111;
12'b0110001101101: data = 6'b111111;
12'b0110001101110: data = 6'b111111;
12'b0110001101111: data = 6'b111111;
12'b0110001110000: data = 6'b111111;
12'b0110001110001: data = 6'b111111;
12'b0110001110010: data = 6'b111111;
12'b0110001110011: data = 6'b111111;
12'b0110001110100: data = 6'b111111;
12'b0110001110101: data = 6'b111111;
12'b0110001110110: data = 6'b111111;
12'b0110001110111: data = 6'b111111;
12'b0110001111000: data = 6'b111111;
12'b0110001111001: data = 6'b111111;
12'b0110001111010: data = 6'b111111;
12'b0110001111011: data = 6'b111111;
12'b0110001111100: data = 6'b111111;
12'b0110001111101: data = 6'b111111;
12'b0110001111110: data = 6'b111111;
12'b0110001111111: data = 6'b111111;
12'b01100010000000: data = 6'b111111;
12'b01100010000001: data = 6'b111111;
12'b01100010000010: data = 6'b111111;
12'b01100010000011: data = 6'b111111;
12'b01100010000100: data = 6'b111111;
12'b01100010000101: data = 6'b111111;
12'b01100010000110: data = 6'b111111;
12'b01100010000111: data = 6'b111111;
12'b01100010001000: data = 6'b111111;
12'b01100010001001: data = 6'b111111;
12'b01100010001010: data = 6'b111111;
12'b01100010001011: data = 6'b010101;
12'b01100010001100: data = 6'b000000;
12'b01100010001101: data = 6'b000000;
12'b01100010001110: data = 6'b101010;
12'b01100010001111: data = 6'b101010;
12'b01100010010000: data = 6'b101010;
12'b01100010010001: data = 6'b101010;
12'b01100010010010: data = 6'b010101;
12'b01100010010011: data = 6'b010101;
12'b01100010010100: data = 6'b010101;
12'b01100010010101: data = 6'b010101;
12'b01100010010110: data = 6'b010101;
12'b01100010010111: data = 6'b010101;
12'b01100010011000: data = 6'b010101;
12'b01100010011001: data = 6'b010101;
12'b01100010011010: data = 6'b010101;
12'b01100010011011: data = 6'b010101;
12'b01100010011100: data = 6'b010101;
12'b01100010011101: data = 6'b010101;
12'b01100010011110: data = 6'b010101;
12'b01100010011111: data = 6'b010101;
12'b01100010100000: data = 6'b010101;
12'b01100010100001: data = 6'b010101;
12'b01100010100010: data = 6'b010101;
12'b01100010100011: data = 6'b010101;
12'b01100010100100: data = 6'b010101;
12'b01100010100101: data = 6'b010101;
12'b01100010100110: data = 6'b010101;
12'b01100010100111: data = 6'b010101;
12'b01100010101000: data = 6'b010101;
12'b01100010101001: data = 6'b010101;
12'b01100010101010: data = 6'b010101;
12'b011001000000: data = 6'b010101;
12'b011001000001: data = 6'b010101;
12'b011001000010: data = 6'b010101;
12'b011001000011: data = 6'b010101;
12'b011001000100: data = 6'b010101;
12'b011001000101: data = 6'b010101;
12'b011001000110: data = 6'b010101;
12'b011001000111: data = 6'b010101;
12'b011001001000: data = 6'b010101;
12'b011001001001: data = 6'b010101;
12'b011001001010: data = 6'b010101;
12'b011001001011: data = 6'b010101;
12'b011001001100: data = 6'b010101;
12'b011001001101: data = 6'b010101;
12'b011001001110: data = 6'b010101;
12'b011001001111: data = 6'b010101;
12'b011001010000: data = 6'b010101;
12'b011001010001: data = 6'b010101;
12'b011001010010: data = 6'b010101;
12'b011001010011: data = 6'b010101;
12'b011001010100: data = 6'b010101;
12'b011001010101: data = 6'b010101;
12'b011001010110: data = 6'b010101;
12'b011001010111: data = 6'b010101;
12'b011001011000: data = 6'b010101;
12'b011001011001: data = 6'b101010;
12'b011001011010: data = 6'b101010;
12'b011001011011: data = 6'b101010;
12'b011001011100: data = 6'b010101;
12'b011001011101: data = 6'b000000;
12'b011001011110: data = 6'b000000;
12'b011001011111: data = 6'b010101;
12'b011001100000: data = 6'b111111;
12'b011001100001: data = 6'b111111;
12'b011001100010: data = 6'b111111;
12'b011001100011: data = 6'b111111;
12'b011001100100: data = 6'b111111;
12'b011001100101: data = 6'b111111;
12'b011001100110: data = 6'b111111;
12'b011001100111: data = 6'b111111;
12'b011001101000: data = 6'b111111;
12'b011001101001: data = 6'b111111;
12'b011001101010: data = 6'b111111;
12'b011001101011: data = 6'b111111;
12'b011001101100: data = 6'b111111;
12'b011001101101: data = 6'b111111;
12'b011001101110: data = 6'b111111;
12'b011001101111: data = 6'b111111;
12'b011001110000: data = 6'b111111;
12'b011001110001: data = 6'b111111;
12'b011001110010: data = 6'b111111;
12'b011001110011: data = 6'b111111;
12'b011001110100: data = 6'b111111;
12'b011001110101: data = 6'b111111;
12'b011001110110: data = 6'b111111;
12'b011001110111: data = 6'b111111;
12'b011001111000: data = 6'b111111;
12'b011001111001: data = 6'b111111;
12'b011001111010: data = 6'b111111;
12'b011001111011: data = 6'b111111;
12'b011001111100: data = 6'b111111;
12'b011001111101: data = 6'b111111;
12'b011001111110: data = 6'b111111;
12'b011001111111: data = 6'b111111;
12'b0110011000000: data = 6'b111111;
12'b0110011000001: data = 6'b111111;
12'b0110011000010: data = 6'b111111;
12'b0110011000011: data = 6'b111111;
12'b0110011000100: data = 6'b111111;
12'b0110011000101: data = 6'b111111;
12'b0110011000110: data = 6'b111111;
12'b0110011000111: data = 6'b111111;
12'b0110011001000: data = 6'b111111;
12'b0110011001001: data = 6'b111111;
12'b0110011001010: data = 6'b111111;
12'b0110011001011: data = 6'b111111;
12'b0110011001100: data = 6'b111111;
12'b0110011001101: data = 6'b111111;
12'b0110011001110: data = 6'b111111;
12'b0110011001111: data = 6'b111111;
12'b0110011010000: data = 6'b111111;
12'b0110011010001: data = 6'b111111;
12'b0110011010010: data = 6'b111111;
12'b0110011010011: data = 6'b111111;
12'b0110011010100: data = 6'b111111;
12'b0110011010101: data = 6'b111111;
12'b0110011010110: data = 6'b111111;
12'b0110011010111: data = 6'b111111;
12'b0110011011000: data = 6'b111111;
12'b0110011011001: data = 6'b111111;
12'b0110011011010: data = 6'b111111;
12'b0110011011011: data = 6'b111111;
12'b0110011011100: data = 6'b111111;
12'b0110011011101: data = 6'b111111;
12'b0110011011110: data = 6'b111111;
12'b0110011011111: data = 6'b111111;
12'b0110011100000: data = 6'b111111;
12'b0110011100001: data = 6'b111111;
12'b0110011100010: data = 6'b111111;
12'b0110011100011: data = 6'b111111;
12'b0110011100100: data = 6'b111111;
12'b0110011100101: data = 6'b111111;
12'b0110011100110: data = 6'b111111;
12'b0110011100111: data = 6'b111111;
12'b0110011101000: data = 6'b111111;
12'b0110011101001: data = 6'b111111;
12'b0110011101010: data = 6'b111111;
12'b0110011101011: data = 6'b111111;
12'b0110011101100: data = 6'b111111;
12'b0110011101101: data = 6'b111111;
12'b0110011101110: data = 6'b111111;
12'b0110011101111: data = 6'b111111;
12'b0110011110000: data = 6'b111111;
12'b0110011110001: data = 6'b111111;
12'b0110011110010: data = 6'b111111;
12'b0110011110011: data = 6'b111111;
12'b0110011110100: data = 6'b111111;
12'b0110011110101: data = 6'b111111;
12'b0110011110110: data = 6'b111111;
12'b0110011110111: data = 6'b111111;
12'b0110011111000: data = 6'b111111;
12'b0110011111001: data = 6'b111111;
12'b0110011111010: data = 6'b111111;
12'b0110011111011: data = 6'b111111;
12'b0110011111100: data = 6'b111111;
12'b0110011111101: data = 6'b111111;
12'b0110011111110: data = 6'b111111;
12'b0110011111111: data = 6'b111111;
12'b01100110000000: data = 6'b111111;
12'b01100110000001: data = 6'b111111;
12'b01100110000010: data = 6'b111111;
12'b01100110000011: data = 6'b111111;
12'b01100110000100: data = 6'b111111;
12'b01100110000101: data = 6'b111111;
12'b01100110000110: data = 6'b111111;
12'b01100110000111: data = 6'b111111;
12'b01100110001000: data = 6'b111111;
12'b01100110001001: data = 6'b111111;
12'b01100110001010: data = 6'b111111;
12'b01100110001011: data = 6'b010101;
12'b01100110001100: data = 6'b000000;
12'b01100110001101: data = 6'b000000;
12'b01100110001110: data = 6'b101010;
12'b01100110001111: data = 6'b101010;
12'b01100110010000: data = 6'b101010;
12'b01100110010001: data = 6'b101010;
12'b01100110010010: data = 6'b010101;
12'b01100110010011: data = 6'b010101;
12'b01100110010100: data = 6'b010101;
12'b01100110010101: data = 6'b010101;
12'b01100110010110: data = 6'b010101;
12'b01100110010111: data = 6'b010101;
12'b01100110011000: data = 6'b010101;
12'b01100110011001: data = 6'b010101;
12'b01100110011010: data = 6'b010101;
12'b01100110011011: data = 6'b010101;
12'b01100110011100: data = 6'b010101;
12'b01100110011101: data = 6'b010101;
12'b01100110011110: data = 6'b010101;
12'b01100110011111: data = 6'b010101;
12'b01100110100000: data = 6'b010101;
12'b01100110100001: data = 6'b010101;
12'b01100110100010: data = 6'b010101;
12'b01100110100011: data = 6'b010101;
12'b01100110100100: data = 6'b010101;
12'b01100110100101: data = 6'b010101;
12'b01100110100110: data = 6'b010101;
12'b01100110100111: data = 6'b010101;
12'b01100110101000: data = 6'b010101;
12'b01100110101001: data = 6'b010101;
12'b01100110101010: data = 6'b010101;
12'b011010000000: data = 6'b010101;
12'b011010000001: data = 6'b010101;
12'b011010000010: data = 6'b010101;
12'b011010000011: data = 6'b010101;
12'b011010000100: data = 6'b010101;
12'b011010000101: data = 6'b010101;
12'b011010000110: data = 6'b010101;
12'b011010000111: data = 6'b010101;
12'b011010001000: data = 6'b010101;
12'b011010001001: data = 6'b010101;
12'b011010001010: data = 6'b010101;
12'b011010001011: data = 6'b010101;
12'b011010001100: data = 6'b010101;
12'b011010001101: data = 6'b010101;
12'b011010001110: data = 6'b010101;
12'b011010001111: data = 6'b010101;
12'b011010010000: data = 6'b010101;
12'b011010010001: data = 6'b010101;
12'b011010010010: data = 6'b010101;
12'b011010010011: data = 6'b010101;
12'b011010010100: data = 6'b010101;
12'b011010010101: data = 6'b010101;
12'b011010010110: data = 6'b010101;
12'b011010010111: data = 6'b010101;
12'b011010011000: data = 6'b010101;
12'b011010011001: data = 6'b101010;
12'b011010011010: data = 6'b101010;
12'b011010011011: data = 6'b101010;
12'b011010011100: data = 6'b010101;
12'b011010011101: data = 6'b000000;
12'b011010011110: data = 6'b000000;
12'b011010011111: data = 6'b010101;
12'b011010100000: data = 6'b101010;
12'b011010100001: data = 6'b101010;
12'b011010100010: data = 6'b111111;
12'b011010100011: data = 6'b111111;
12'b011010100100: data = 6'b111111;
12'b011010100101: data = 6'b111111;
12'b011010100110: data = 6'b111111;
12'b011010100111: data = 6'b111111;
12'b011010101000: data = 6'b111111;
12'b011010101001: data = 6'b111111;
12'b011010101010: data = 6'b111111;
12'b011010101011: data = 6'b111111;
12'b011010101100: data = 6'b111111;
12'b011010101101: data = 6'b111111;
12'b011010101110: data = 6'b111111;
12'b011010101111: data = 6'b111111;
12'b011010110000: data = 6'b111111;
12'b011010110001: data = 6'b111111;
12'b011010110010: data = 6'b111111;
12'b011010110011: data = 6'b111111;
12'b011010110100: data = 6'b111111;
12'b011010110101: data = 6'b111111;
12'b011010110110: data = 6'b111111;
12'b011010110111: data = 6'b111111;
12'b011010111000: data = 6'b111111;
12'b011010111001: data = 6'b111111;
12'b011010111010: data = 6'b111111;
12'b011010111011: data = 6'b111111;
12'b011010111100: data = 6'b111111;
12'b011010111101: data = 6'b111111;
12'b011010111110: data = 6'b111111;
12'b011010111111: data = 6'b111111;
12'b0110101000000: data = 6'b111111;
12'b0110101000001: data = 6'b111111;
12'b0110101000010: data = 6'b111111;
12'b0110101000011: data = 6'b111111;
12'b0110101000100: data = 6'b111111;
12'b0110101000101: data = 6'b111111;
12'b0110101000110: data = 6'b111111;
12'b0110101000111: data = 6'b111111;
12'b0110101001000: data = 6'b111111;
12'b0110101001001: data = 6'b111111;
12'b0110101001010: data = 6'b111111;
12'b0110101001011: data = 6'b111111;
12'b0110101001100: data = 6'b111111;
12'b0110101001101: data = 6'b111111;
12'b0110101001110: data = 6'b111111;
12'b0110101001111: data = 6'b111111;
12'b0110101010000: data = 6'b111111;
12'b0110101010001: data = 6'b111111;
12'b0110101010010: data = 6'b111111;
12'b0110101010011: data = 6'b111111;
12'b0110101010100: data = 6'b111111;
12'b0110101010101: data = 6'b111111;
12'b0110101010110: data = 6'b111111;
12'b0110101010111: data = 6'b111111;
12'b0110101011000: data = 6'b111111;
12'b0110101011001: data = 6'b111111;
12'b0110101011010: data = 6'b111111;
12'b0110101011011: data = 6'b111111;
12'b0110101011100: data = 6'b111111;
12'b0110101011101: data = 6'b111111;
12'b0110101011110: data = 6'b111111;
12'b0110101011111: data = 6'b111111;
12'b0110101100000: data = 6'b111111;
12'b0110101100001: data = 6'b111111;
12'b0110101100010: data = 6'b111111;
12'b0110101100011: data = 6'b111111;
12'b0110101100100: data = 6'b111111;
12'b0110101100101: data = 6'b111111;
12'b0110101100110: data = 6'b111111;
12'b0110101100111: data = 6'b111111;
12'b0110101101000: data = 6'b111111;
12'b0110101101001: data = 6'b111111;
12'b0110101101010: data = 6'b111111;
12'b0110101101011: data = 6'b111111;
12'b0110101101100: data = 6'b111111;
12'b0110101101101: data = 6'b111111;
12'b0110101101110: data = 6'b111111;
12'b0110101101111: data = 6'b111111;
12'b0110101110000: data = 6'b111111;
12'b0110101110001: data = 6'b111111;
12'b0110101110010: data = 6'b111111;
12'b0110101110011: data = 6'b111111;
12'b0110101110100: data = 6'b111111;
12'b0110101110101: data = 6'b111111;
12'b0110101110110: data = 6'b111111;
12'b0110101110111: data = 6'b111111;
12'b0110101111000: data = 6'b111111;
12'b0110101111001: data = 6'b111111;
12'b0110101111010: data = 6'b111111;
12'b0110101111011: data = 6'b111111;
12'b0110101111100: data = 6'b111111;
12'b0110101111101: data = 6'b111111;
12'b0110101111110: data = 6'b111111;
12'b0110101111111: data = 6'b111111;
12'b01101010000000: data = 6'b111111;
12'b01101010000001: data = 6'b111111;
12'b01101010000010: data = 6'b111111;
12'b01101010000011: data = 6'b111111;
12'b01101010000100: data = 6'b111111;
12'b01101010000101: data = 6'b111111;
12'b01101010000110: data = 6'b111111;
12'b01101010000111: data = 6'b111111;
12'b01101010001000: data = 6'b111111;
12'b01101010001001: data = 6'b101010;
12'b01101010001010: data = 6'b101010;
12'b01101010001011: data = 6'b010101;
12'b01101010001100: data = 6'b000000;
12'b01101010001101: data = 6'b000000;
12'b01101010001110: data = 6'b101010;
12'b01101010001111: data = 6'b101010;
12'b01101010010000: data = 6'b101010;
12'b01101010010001: data = 6'b101010;
12'b01101010010010: data = 6'b010101;
12'b01101010010011: data = 6'b010101;
12'b01101010010100: data = 6'b010101;
12'b01101010010101: data = 6'b010101;
12'b01101010010110: data = 6'b010101;
12'b01101010010111: data = 6'b010101;
12'b01101010011000: data = 6'b010101;
12'b01101010011001: data = 6'b010101;
12'b01101010011010: data = 6'b010101;
12'b01101010011011: data = 6'b010101;
12'b01101010011100: data = 6'b010101;
12'b01101010011101: data = 6'b010101;
12'b01101010011110: data = 6'b010101;
12'b01101010011111: data = 6'b010101;
12'b01101010100000: data = 6'b010101;
12'b01101010100001: data = 6'b010101;
12'b01101010100010: data = 6'b010101;
12'b01101010100011: data = 6'b010101;
12'b01101010100100: data = 6'b010101;
12'b01101010100101: data = 6'b010101;
12'b01101010100110: data = 6'b010101;
12'b01101010100111: data = 6'b010101;
12'b01101010101000: data = 6'b010101;
12'b01101010101001: data = 6'b010101;
12'b01101010101010: data = 6'b010101;
12'b011011000000: data = 6'b010101;
12'b011011000001: data = 6'b010101;
12'b011011000010: data = 6'b010101;
12'b011011000011: data = 6'b010101;
12'b011011000100: data = 6'b010101;
12'b011011000101: data = 6'b010101;
12'b011011000110: data = 6'b010101;
12'b011011000111: data = 6'b010101;
12'b011011001000: data = 6'b010101;
12'b011011001001: data = 6'b010101;
12'b011011001010: data = 6'b010101;
12'b011011001011: data = 6'b010101;
12'b011011001100: data = 6'b010101;
12'b011011001101: data = 6'b010101;
12'b011011001110: data = 6'b010101;
12'b011011001111: data = 6'b010101;
12'b011011010000: data = 6'b010101;
12'b011011010001: data = 6'b010101;
12'b011011010010: data = 6'b010101;
12'b011011010011: data = 6'b010101;
12'b011011010100: data = 6'b010101;
12'b011011010101: data = 6'b010101;
12'b011011010110: data = 6'b010101;
12'b011011010111: data = 6'b010101;
12'b011011011000: data = 6'b010101;
12'b011011011001: data = 6'b101010;
12'b011011011010: data = 6'b101010;
12'b011011011011: data = 6'b101010;
12'b011011011100: data = 6'b010101;
12'b011011011101: data = 6'b000000;
12'b011011011110: data = 6'b000000;
12'b011011011111: data = 6'b000000;
12'b011011100000: data = 6'b010101;
12'b011011100001: data = 6'b010101;
12'b011011100010: data = 6'b101010;
12'b011011100011: data = 6'b111111;
12'b011011100100: data = 6'b111111;
12'b011011100101: data = 6'b111111;
12'b011011100110: data = 6'b111111;
12'b011011100111: data = 6'b111111;
12'b011011101000: data = 6'b111111;
12'b011011101001: data = 6'b111111;
12'b011011101010: data = 6'b111111;
12'b011011101011: data = 6'b111111;
12'b011011101100: data = 6'b111111;
12'b011011101101: data = 6'b111111;
12'b011011101110: data = 6'b111111;
12'b011011101111: data = 6'b111111;
12'b011011110000: data = 6'b111111;
12'b011011110001: data = 6'b111111;
12'b011011110010: data = 6'b111111;
12'b011011110011: data = 6'b111111;
12'b011011110100: data = 6'b111111;
12'b011011110101: data = 6'b111111;
12'b011011110110: data = 6'b111111;
12'b011011110111: data = 6'b111111;
12'b011011111000: data = 6'b111111;
12'b011011111001: data = 6'b111111;
12'b011011111010: data = 6'b111111;
12'b011011111011: data = 6'b111111;
12'b011011111100: data = 6'b111111;
12'b011011111101: data = 6'b111111;
12'b011011111110: data = 6'b111111;
12'b011011111111: data = 6'b111111;
12'b0110111000000: data = 6'b111111;
12'b0110111000001: data = 6'b111111;
12'b0110111000010: data = 6'b111111;
12'b0110111000011: data = 6'b111111;
12'b0110111000100: data = 6'b111111;
12'b0110111000101: data = 6'b111111;
12'b0110111000110: data = 6'b111111;
12'b0110111000111: data = 6'b111111;
12'b0110111001000: data = 6'b111111;
12'b0110111001001: data = 6'b111111;
12'b0110111001010: data = 6'b111111;
12'b0110111001011: data = 6'b111111;
12'b0110111001100: data = 6'b111111;
12'b0110111001101: data = 6'b111111;
12'b0110111001110: data = 6'b111111;
12'b0110111001111: data = 6'b111111;
12'b0110111010000: data = 6'b111111;
12'b0110111010001: data = 6'b111111;
12'b0110111010010: data = 6'b111111;
12'b0110111010011: data = 6'b111111;
12'b0110111010100: data = 6'b111111;
12'b0110111010101: data = 6'b111111;
12'b0110111010110: data = 6'b111111;
12'b0110111010111: data = 6'b111111;
12'b0110111011000: data = 6'b111111;
12'b0110111011001: data = 6'b111111;
12'b0110111011010: data = 6'b111111;
12'b0110111011011: data = 6'b111111;
12'b0110111011100: data = 6'b111111;
12'b0110111011101: data = 6'b111111;
12'b0110111011110: data = 6'b111111;
12'b0110111011111: data = 6'b111111;
12'b0110111100000: data = 6'b111111;
12'b0110111100001: data = 6'b111111;
12'b0110111100010: data = 6'b111111;
12'b0110111100011: data = 6'b111111;
12'b0110111100100: data = 6'b111111;
12'b0110111100101: data = 6'b111111;
12'b0110111100110: data = 6'b111111;
12'b0110111100111: data = 6'b111111;
12'b0110111101000: data = 6'b111111;
12'b0110111101001: data = 6'b111111;
12'b0110111101010: data = 6'b111111;
12'b0110111101011: data = 6'b111111;
12'b0110111101100: data = 6'b111111;
12'b0110111101101: data = 6'b111111;
12'b0110111101110: data = 6'b111111;
12'b0110111101111: data = 6'b111111;
12'b0110111110000: data = 6'b111111;
12'b0110111110001: data = 6'b111111;
12'b0110111110010: data = 6'b111111;
12'b0110111110011: data = 6'b111111;
12'b0110111110100: data = 6'b111111;
12'b0110111110101: data = 6'b111111;
12'b0110111110110: data = 6'b111111;
12'b0110111110111: data = 6'b111111;
12'b0110111111000: data = 6'b111111;
12'b0110111111001: data = 6'b111111;
12'b0110111111010: data = 6'b111111;
12'b0110111111011: data = 6'b111111;
12'b0110111111100: data = 6'b111111;
12'b0110111111101: data = 6'b111111;
12'b0110111111110: data = 6'b111111;
12'b0110111111111: data = 6'b111111;
12'b01101110000000: data = 6'b111111;
12'b01101110000001: data = 6'b111111;
12'b01101110000010: data = 6'b111111;
12'b01101110000011: data = 6'b111111;
12'b01101110000100: data = 6'b111111;
12'b01101110000101: data = 6'b111111;
12'b01101110000110: data = 6'b111111;
12'b01101110000111: data = 6'b111111;
12'b01101110001000: data = 6'b111111;
12'b01101110001001: data = 6'b101010;
12'b01101110001010: data = 6'b101010;
12'b01101110001011: data = 6'b010101;
12'b01101110001100: data = 6'b000000;
12'b01101110001101: data = 6'b000000;
12'b01101110001110: data = 6'b101010;
12'b01101110001111: data = 6'b101010;
12'b01101110010000: data = 6'b101010;
12'b01101110010001: data = 6'b101010;
12'b01101110010010: data = 6'b010101;
12'b01101110010011: data = 6'b010101;
12'b01101110010100: data = 6'b010101;
12'b01101110010101: data = 6'b010101;
12'b01101110010110: data = 6'b010101;
12'b01101110010111: data = 6'b010101;
12'b01101110011000: data = 6'b010101;
12'b01101110011001: data = 6'b010101;
12'b01101110011010: data = 6'b010101;
12'b01101110011011: data = 6'b010101;
12'b01101110011100: data = 6'b010101;
12'b01101110011101: data = 6'b010101;
12'b01101110011110: data = 6'b010101;
12'b01101110011111: data = 6'b010101;
12'b01101110100000: data = 6'b010101;
12'b01101110100001: data = 6'b010101;
12'b01101110100010: data = 6'b010101;
12'b01101110100011: data = 6'b010101;
12'b01101110100100: data = 6'b010101;
12'b01101110100101: data = 6'b010101;
12'b01101110100110: data = 6'b010101;
12'b01101110100111: data = 6'b010101;
12'b01101110101000: data = 6'b010101;
12'b01101110101001: data = 6'b010101;
12'b01101110101010: data = 6'b010101;
12'b011100000000: data = 6'b010101;
12'b011100000001: data = 6'b010101;
12'b011100000010: data = 6'b010101;
12'b011100000011: data = 6'b010101;
12'b011100000100: data = 6'b010101;
12'b011100000101: data = 6'b010101;
12'b011100000110: data = 6'b010101;
12'b011100000111: data = 6'b010101;
12'b011100001000: data = 6'b010101;
12'b011100001001: data = 6'b010101;
12'b011100001010: data = 6'b010101;
12'b011100001011: data = 6'b010101;
12'b011100001100: data = 6'b010101;
12'b011100001101: data = 6'b010101;
12'b011100001110: data = 6'b010101;
12'b011100001111: data = 6'b010101;
12'b011100010000: data = 6'b010101;
12'b011100010001: data = 6'b010101;
12'b011100010010: data = 6'b010101;
12'b011100010011: data = 6'b010101;
12'b011100010100: data = 6'b010101;
12'b011100010101: data = 6'b010101;
12'b011100010110: data = 6'b010101;
12'b011100010111: data = 6'b010101;
12'b011100011000: data = 6'b010101;
12'b011100011001: data = 6'b101010;
12'b011100011010: data = 6'b101010;
12'b011100011011: data = 6'b101010;
12'b011100011100: data = 6'b010101;
12'b011100011101: data = 6'b000000;
12'b011100011110: data = 6'b000000;
12'b011100011111: data = 6'b000000;
12'b011100100000: data = 6'b010101;
12'b011100100001: data = 6'b010101;
12'b011100100010: data = 6'b101010;
12'b011100100011: data = 6'b111111;
12'b011100100100: data = 6'b111111;
12'b011100100101: data = 6'b111111;
12'b011100100110: data = 6'b111111;
12'b011100100111: data = 6'b111111;
12'b011100101000: data = 6'b111111;
12'b011100101001: data = 6'b111111;
12'b011100101010: data = 6'b111111;
12'b011100101011: data = 6'b111111;
12'b011100101100: data = 6'b111111;
12'b011100101101: data = 6'b111111;
12'b011100101110: data = 6'b111111;
12'b011100101111: data = 6'b111111;
12'b011100110000: data = 6'b111111;
12'b011100110001: data = 6'b111111;
12'b011100110010: data = 6'b111111;
12'b011100110011: data = 6'b111111;
12'b011100110100: data = 6'b111111;
12'b011100110101: data = 6'b111111;
12'b011100110110: data = 6'b111111;
12'b011100110111: data = 6'b111111;
12'b011100111000: data = 6'b111111;
12'b011100111001: data = 6'b111111;
12'b011100111010: data = 6'b111111;
12'b011100111011: data = 6'b111111;
12'b011100111100: data = 6'b111111;
12'b011100111101: data = 6'b111111;
12'b011100111110: data = 6'b111111;
12'b011100111111: data = 6'b111111;
12'b0111001000000: data = 6'b111111;
12'b0111001000001: data = 6'b111111;
12'b0111001000010: data = 6'b111111;
12'b0111001000011: data = 6'b111111;
12'b0111001000100: data = 6'b111111;
12'b0111001000101: data = 6'b111111;
12'b0111001000110: data = 6'b111111;
12'b0111001000111: data = 6'b111111;
12'b0111001001000: data = 6'b111111;
12'b0111001001001: data = 6'b111111;
12'b0111001001010: data = 6'b111111;
12'b0111001001011: data = 6'b111111;
12'b0111001001100: data = 6'b111111;
12'b0111001001101: data = 6'b111111;
12'b0111001001110: data = 6'b111111;
12'b0111001001111: data = 6'b111111;
12'b0111001010000: data = 6'b111111;
12'b0111001010001: data = 6'b111111;
12'b0111001010010: data = 6'b111111;
12'b0111001010011: data = 6'b111111;
12'b0111001010100: data = 6'b111111;
12'b0111001010101: data = 6'b111111;
12'b0111001010110: data = 6'b111111;
12'b0111001010111: data = 6'b111111;
12'b0111001011000: data = 6'b111111;
12'b0111001011001: data = 6'b111111;
12'b0111001011010: data = 6'b111111;
12'b0111001011011: data = 6'b111111;
12'b0111001011100: data = 6'b111111;
12'b0111001011101: data = 6'b111111;
12'b0111001011110: data = 6'b111111;
12'b0111001011111: data = 6'b111111;
12'b0111001100000: data = 6'b111111;
12'b0111001100001: data = 6'b111111;
12'b0111001100010: data = 6'b111111;
12'b0111001100011: data = 6'b111111;
12'b0111001100100: data = 6'b111111;
12'b0111001100101: data = 6'b111111;
12'b0111001100110: data = 6'b111111;
12'b0111001100111: data = 6'b111111;
12'b0111001101000: data = 6'b111111;
12'b0111001101001: data = 6'b111111;
12'b0111001101010: data = 6'b111111;
12'b0111001101011: data = 6'b111111;
12'b0111001101100: data = 6'b111111;
12'b0111001101101: data = 6'b111111;
12'b0111001101110: data = 6'b111111;
12'b0111001101111: data = 6'b111111;
12'b0111001110000: data = 6'b111111;
12'b0111001110001: data = 6'b111111;
12'b0111001110010: data = 6'b111111;
12'b0111001110011: data = 6'b111111;
12'b0111001110100: data = 6'b111111;
12'b0111001110101: data = 6'b111111;
12'b0111001110110: data = 6'b111111;
12'b0111001110111: data = 6'b111111;
12'b0111001111000: data = 6'b111111;
12'b0111001111001: data = 6'b111111;
12'b0111001111010: data = 6'b111111;
12'b0111001111011: data = 6'b111111;
12'b0111001111100: data = 6'b111111;
12'b0111001111101: data = 6'b111111;
12'b0111001111110: data = 6'b111111;
12'b0111001111111: data = 6'b111111;
12'b01110010000000: data = 6'b111111;
12'b01110010000001: data = 6'b111111;
12'b01110010000010: data = 6'b111111;
12'b01110010000011: data = 6'b111111;
12'b01110010000100: data = 6'b111111;
12'b01110010000101: data = 6'b111111;
12'b01110010000110: data = 6'b111111;
12'b01110010000111: data = 6'b111111;
12'b01110010001000: data = 6'b111111;
12'b01110010001001: data = 6'b101010;
12'b01110010001010: data = 6'b101010;
12'b01110010001011: data = 6'b010101;
12'b01110010001100: data = 6'b000000;
12'b01110010001101: data = 6'b000000;
12'b01110010001110: data = 6'b101010;
12'b01110010001111: data = 6'b101010;
12'b01110010010000: data = 6'b101010;
12'b01110010010001: data = 6'b101010;
12'b01110010010010: data = 6'b010101;
12'b01110010010011: data = 6'b010101;
12'b01110010010100: data = 6'b010101;
12'b01110010010101: data = 6'b010101;
12'b01110010010110: data = 6'b010101;
12'b01110010010111: data = 6'b010101;
12'b01110010011000: data = 6'b010101;
12'b01110010011001: data = 6'b010101;
12'b01110010011010: data = 6'b010101;
12'b01110010011011: data = 6'b010101;
12'b01110010011100: data = 6'b010101;
12'b01110010011101: data = 6'b010101;
12'b01110010011110: data = 6'b010101;
12'b01110010011111: data = 6'b010101;
12'b01110010100000: data = 6'b010101;
12'b01110010100001: data = 6'b010101;
12'b01110010100010: data = 6'b010101;
12'b01110010100011: data = 6'b010101;
12'b01110010100100: data = 6'b010101;
12'b01110010100101: data = 6'b010101;
12'b01110010100110: data = 6'b010101;
12'b01110010100111: data = 6'b010101;
12'b01110010101000: data = 6'b010101;
12'b01110010101001: data = 6'b010101;
12'b01110010101010: data = 6'b010101;
12'b011101000000: data = 6'b010101;
12'b011101000001: data = 6'b010101;
12'b011101000010: data = 6'b010101;
12'b011101000011: data = 6'b010101;
12'b011101000100: data = 6'b010101;
12'b011101000101: data = 6'b010101;
12'b011101000110: data = 6'b010101;
12'b011101000111: data = 6'b010101;
12'b011101001000: data = 6'b010101;
12'b011101001001: data = 6'b010101;
12'b011101001010: data = 6'b010101;
12'b011101001011: data = 6'b010101;
12'b011101001100: data = 6'b010101;
12'b011101001101: data = 6'b010101;
12'b011101001110: data = 6'b010101;
12'b011101001111: data = 6'b010101;
12'b011101010000: data = 6'b010101;
12'b011101010001: data = 6'b010101;
12'b011101010010: data = 6'b010101;
12'b011101010011: data = 6'b010101;
12'b011101010100: data = 6'b010101;
12'b011101010101: data = 6'b010101;
12'b011101010110: data = 6'b010101;
12'b011101010111: data = 6'b010101;
12'b011101011000: data = 6'b010101;
12'b011101011001: data = 6'b101010;
12'b011101011010: data = 6'b101010;
12'b011101011011: data = 6'b101010;
12'b011101011100: data = 6'b101010;
12'b011101011101: data = 6'b010101;
12'b011101011110: data = 6'b010101;
12'b011101011111: data = 6'b010101;
12'b011101100000: data = 6'b010101;
12'b011101100001: data = 6'b010101;
12'b011101100010: data = 6'b101010;
12'b011101100011: data = 6'b101010;
12'b011101100100: data = 6'b101010;
12'b011101100101: data = 6'b101010;
12'b011101100110: data = 6'b101010;
12'b011101100111: data = 6'b010101;
12'b011101101000: data = 6'b010101;
12'b011101101001: data = 6'b010101;
12'b011101101010: data = 6'b010101;
12'b011101101011: data = 6'b010101;
12'b011101101100: data = 6'b010101;
12'b011101101101: data = 6'b010101;
12'b011101101110: data = 6'b010101;
12'b011101101111: data = 6'b010101;
12'b011101110000: data = 6'b010101;
12'b011101110001: data = 6'b010101;
12'b011101110010: data = 6'b010101;
12'b011101110011: data = 6'b010101;
12'b011101110100: data = 6'b010101;
12'b011101110101: data = 6'b010101;
12'b011101110110: data = 6'b010101;
12'b011101110111: data = 6'b010101;
12'b011101111000: data = 6'b010101;
12'b011101111001: data = 6'b010101;
12'b011101111010: data = 6'b010101;
12'b011101111011: data = 6'b010101;
12'b011101111100: data = 6'b010101;
12'b011101111101: data = 6'b010101;
12'b011101111110: data = 6'b010101;
12'b011101111111: data = 6'b010101;
12'b0111011000000: data = 6'b010101;
12'b0111011000001: data = 6'b010101;
12'b0111011000010: data = 6'b010101;
12'b0111011000011: data = 6'b010101;
12'b0111011000100: data = 6'b010101;
12'b0111011000101: data = 6'b010101;
12'b0111011000110: data = 6'b010101;
12'b0111011000111: data = 6'b010101;
12'b0111011001000: data = 6'b010101;
12'b0111011001001: data = 6'b010101;
12'b0111011001010: data = 6'b010101;
12'b0111011001011: data = 6'b010101;
12'b0111011001100: data = 6'b010101;
12'b0111011001101: data = 6'b010101;
12'b0111011001110: data = 6'b010101;
12'b0111011001111: data = 6'b010101;
12'b0111011010000: data = 6'b010101;
12'b0111011010001: data = 6'b010101;
12'b0111011010010: data = 6'b010101;
12'b0111011010011: data = 6'b010101;
12'b0111011010100: data = 6'b010101;
12'b0111011010101: data = 6'b010101;
12'b0111011010110: data = 6'b010101;
12'b0111011010111: data = 6'b010101;
12'b0111011011000: data = 6'b010101;
12'b0111011011001: data = 6'b010101;
12'b0111011011010: data = 6'b010101;
12'b0111011011011: data = 6'b010101;
12'b0111011011100: data = 6'b010101;
12'b0111011011101: data = 6'b010101;
12'b0111011011110: data = 6'b010101;
12'b0111011011111: data = 6'b010101;
12'b0111011100000: data = 6'b010101;
12'b0111011100001: data = 6'b010101;
12'b0111011100010: data = 6'b010101;
12'b0111011100011: data = 6'b010101;
12'b0111011100100: data = 6'b010101;
12'b0111011100101: data = 6'b010101;
12'b0111011100110: data = 6'b010101;
12'b0111011100111: data = 6'b010101;
12'b0111011101000: data = 6'b010101;
12'b0111011101001: data = 6'b010101;
12'b0111011101010: data = 6'b010101;
12'b0111011101011: data = 6'b010101;
12'b0111011101100: data = 6'b010101;
12'b0111011101101: data = 6'b010101;
12'b0111011101110: data = 6'b010101;
12'b0111011101111: data = 6'b010101;
12'b0111011110000: data = 6'b010101;
12'b0111011110001: data = 6'b010101;
12'b0111011110010: data = 6'b010101;
12'b0111011110011: data = 6'b010101;
12'b0111011110100: data = 6'b010101;
12'b0111011110101: data = 6'b010101;
12'b0111011110110: data = 6'b010101;
12'b0111011110111: data = 6'b010101;
12'b0111011111000: data = 6'b010101;
12'b0111011111001: data = 6'b010101;
12'b0111011111010: data = 6'b010101;
12'b0111011111011: data = 6'b010101;
12'b0111011111100: data = 6'b010101;
12'b0111011111101: data = 6'b010101;
12'b0111011111110: data = 6'b010101;
12'b0111011111111: data = 6'b010101;
12'b01110110000000: data = 6'b010101;
12'b01110110000001: data = 6'b010101;
12'b01110110000010: data = 6'b010101;
12'b01110110000011: data = 6'b010101;
12'b01110110000100: data = 6'b101010;
12'b01110110000101: data = 6'b101010;
12'b01110110000110: data = 6'b101010;
12'b01110110000111: data = 6'b101010;
12'b01110110001000: data = 6'b101010;
12'b01110110001001: data = 6'b101010;
12'b01110110001010: data = 6'b101010;
12'b01110110001011: data = 6'b101001;
12'b01110110001100: data = 6'b101001;
12'b01110110001101: data = 6'b101001;
12'b01110110001110: data = 6'b101010;
12'b01110110001111: data = 6'b101010;
12'b01110110010000: data = 6'b101010;
12'b01110110010001: data = 6'b101010;
12'b01110110010010: data = 6'b010101;
12'b01110110010011: data = 6'b010101;
12'b01110110010100: data = 6'b010101;
12'b01110110010101: data = 6'b010101;
12'b01110110010110: data = 6'b010101;
12'b01110110010111: data = 6'b010101;
12'b01110110011000: data = 6'b010101;
12'b01110110011001: data = 6'b010101;
12'b01110110011010: data = 6'b010101;
12'b01110110011011: data = 6'b010101;
12'b01110110011100: data = 6'b010101;
12'b01110110011101: data = 6'b010101;
12'b01110110011110: data = 6'b010101;
12'b01110110011111: data = 6'b010101;
12'b01110110100000: data = 6'b010101;
12'b01110110100001: data = 6'b010101;
12'b01110110100010: data = 6'b010101;
12'b01110110100011: data = 6'b010101;
12'b01110110100100: data = 6'b010101;
12'b01110110100101: data = 6'b010101;
12'b01110110100110: data = 6'b010101;
12'b01110110100111: data = 6'b010101;
12'b01110110101000: data = 6'b010101;
12'b01110110101001: data = 6'b010101;
12'b01110110101010: data = 6'b010101;
12'b011110000000: data = 6'b010101;
12'b011110000001: data = 6'b010101;
12'b011110000010: data = 6'b010101;
12'b011110000011: data = 6'b010101;
12'b011110000100: data = 6'b010101;
12'b011110000101: data = 6'b010101;
12'b011110000110: data = 6'b010101;
12'b011110000111: data = 6'b010101;
12'b011110001000: data = 6'b010101;
12'b011110001001: data = 6'b010101;
12'b011110001010: data = 6'b010101;
12'b011110001011: data = 6'b010101;
12'b011110001100: data = 6'b010101;
12'b011110001101: data = 6'b010101;
12'b011110001110: data = 6'b010101;
12'b011110001111: data = 6'b010101;
12'b011110010000: data = 6'b010101;
12'b011110010001: data = 6'b010101;
12'b011110010010: data = 6'b010101;
12'b011110010011: data = 6'b010101;
12'b011110010100: data = 6'b010101;
12'b011110010101: data = 6'b010101;
12'b011110010110: data = 6'b010101;
12'b011110010111: data = 6'b010101;
12'b011110011000: data = 6'b010101;
12'b011110011001: data = 6'b101010;
12'b011110011010: data = 6'b101010;
12'b011110011011: data = 6'b101010;
12'b011110011100: data = 6'b101010;
12'b011110011101: data = 6'b101010;
12'b011110011110: data = 6'b101010;
12'b011110011111: data = 6'b101010;
12'b011110100000: data = 6'b010101;
12'b011110100001: data = 6'b010101;
12'b011110100010: data = 6'b010101;
12'b011110100011: data = 6'b010101;
12'b011110100100: data = 6'b010101;
12'b011110100101: data = 6'b010101;
12'b011110100110: data = 6'b010101;
12'b011110100111: data = 6'b000000;
12'b011110101000: data = 6'b000000;
12'b011110101001: data = 6'b000000;
12'b011110101010: data = 6'b000000;
12'b011110101011: data = 6'b000000;
12'b011110101100: data = 6'b000000;
12'b011110101101: data = 6'b000000;
12'b011110101110: data = 6'b000000;
12'b011110101111: data = 6'b000000;
12'b011110110000: data = 6'b000000;
12'b011110110001: data = 6'b000000;
12'b011110110010: data = 6'b000000;
12'b011110110011: data = 6'b000000;
12'b011110110100: data = 6'b000000;
12'b011110110101: data = 6'b000000;
12'b011110110110: data = 6'b000000;
12'b011110110111: data = 6'b000000;
12'b011110111000: data = 6'b000000;
12'b011110111001: data = 6'b000000;
12'b011110111010: data = 6'b000000;
12'b011110111011: data = 6'b000000;
12'b011110111100: data = 6'b000000;
12'b011110111101: data = 6'b000000;
12'b011110111110: data = 6'b000000;
12'b011110111111: data = 6'b000000;
12'b0111101000000: data = 6'b000000;
12'b0111101000001: data = 6'b000000;
12'b0111101000010: data = 6'b000000;
12'b0111101000011: data = 6'b000000;
12'b0111101000100: data = 6'b000000;
12'b0111101000101: data = 6'b000000;
12'b0111101000110: data = 6'b000000;
12'b0111101000111: data = 6'b000000;
12'b0111101001000: data = 6'b000000;
12'b0111101001001: data = 6'b000000;
12'b0111101001010: data = 6'b000000;
12'b0111101001011: data = 6'b000000;
12'b0111101001100: data = 6'b000000;
12'b0111101001101: data = 6'b000000;
12'b0111101001110: data = 6'b000000;
12'b0111101001111: data = 6'b000000;
12'b0111101010000: data = 6'b000000;
12'b0111101010001: data = 6'b000000;
12'b0111101010010: data = 6'b000000;
12'b0111101010011: data = 6'b000000;
12'b0111101010100: data = 6'b000000;
12'b0111101010101: data = 6'b000000;
12'b0111101010110: data = 6'b000000;
12'b0111101010111: data = 6'b000000;
12'b0111101011000: data = 6'b000000;
12'b0111101011001: data = 6'b000000;
12'b0111101011010: data = 6'b000000;
12'b0111101011011: data = 6'b000000;
12'b0111101011100: data = 6'b000000;
12'b0111101011101: data = 6'b000000;
12'b0111101011110: data = 6'b000000;
12'b0111101011111: data = 6'b000000;
12'b0111101100000: data = 6'b000000;
12'b0111101100001: data = 6'b000000;
12'b0111101100010: data = 6'b000000;
12'b0111101100011: data = 6'b000000;
12'b0111101100100: data = 6'b000000;
12'b0111101100101: data = 6'b000000;
12'b0111101100110: data = 6'b000000;
12'b0111101100111: data = 6'b000000;
12'b0111101101000: data = 6'b000000;
12'b0111101101001: data = 6'b000000;
12'b0111101101010: data = 6'b000000;
12'b0111101101011: data = 6'b000000;
12'b0111101101100: data = 6'b000000;
12'b0111101101101: data = 6'b000000;
12'b0111101101110: data = 6'b000000;
12'b0111101101111: data = 6'b000000;
12'b0111101110000: data = 6'b000000;
12'b0111101110001: data = 6'b000000;
12'b0111101110010: data = 6'b000000;
12'b0111101110011: data = 6'b000000;
12'b0111101110100: data = 6'b000000;
12'b0111101110101: data = 6'b000000;
12'b0111101110110: data = 6'b000000;
12'b0111101110111: data = 6'b000000;
12'b0111101111000: data = 6'b000000;
12'b0111101111001: data = 6'b000000;
12'b0111101111010: data = 6'b000000;
12'b0111101111011: data = 6'b000000;
12'b0111101111100: data = 6'b000000;
12'b0111101111101: data = 6'b000000;
12'b0111101111110: data = 6'b000000;
12'b0111101111111: data = 6'b000000;
12'b01111010000000: data = 6'b000000;
12'b01111010000001: data = 6'b000000;
12'b01111010000010: data = 6'b000000;
12'b01111010000011: data = 6'b000000;
12'b01111010000100: data = 6'b000000;
12'b01111010000101: data = 6'b000000;
12'b01111010000110: data = 6'b010101;
12'b01111010000111: data = 6'b010101;
12'b01111010001000: data = 6'b010101;
12'b01111010001001: data = 6'b010101;
12'b01111010001010: data = 6'b010101;
12'b01111010001011: data = 6'b101010;
12'b01111010001100: data = 6'b111111;
12'b01111010001101: data = 6'b111111;
12'b01111010001110: data = 6'b101010;
12'b01111010001111: data = 6'b101010;
12'b01111010010000: data = 6'b101010;
12'b01111010010001: data = 6'b101010;
12'b01111010010010: data = 6'b010101;
12'b01111010010011: data = 6'b010101;
12'b01111010010100: data = 6'b010101;
12'b01111010010101: data = 6'b010101;
12'b01111010010110: data = 6'b010101;
12'b01111010010111: data = 6'b010101;
12'b01111010011000: data = 6'b010101;
12'b01111010011001: data = 6'b010101;
12'b01111010011010: data = 6'b010101;
12'b01111010011011: data = 6'b010101;
12'b01111010011100: data = 6'b010101;
12'b01111010011101: data = 6'b010101;
12'b01111010011110: data = 6'b010101;
12'b01111010011111: data = 6'b010101;
12'b01111010100000: data = 6'b010101;
12'b01111010100001: data = 6'b010101;
12'b01111010100010: data = 6'b010101;
12'b01111010100011: data = 6'b010101;
12'b01111010100100: data = 6'b010101;
12'b01111010100101: data = 6'b010101;
12'b01111010100110: data = 6'b010101;
12'b01111010100111: data = 6'b010101;
12'b01111010101000: data = 6'b010101;
12'b01111010101001: data = 6'b010101;
12'b01111010101010: data = 6'b010101;
12'b011111000000: data = 6'b010101;
12'b011111000001: data = 6'b010101;
12'b011111000010: data = 6'b010101;
12'b011111000011: data = 6'b010101;
12'b011111000100: data = 6'b010101;
12'b011111000101: data = 6'b010101;
12'b011111000110: data = 6'b010101;
12'b011111000111: data = 6'b010101;
12'b011111001000: data = 6'b010101;
12'b011111001001: data = 6'b010101;
12'b011111001010: data = 6'b010101;
12'b011111001011: data = 6'b010101;
12'b011111001100: data = 6'b010101;
12'b011111001101: data = 6'b010101;
12'b011111001110: data = 6'b010101;
12'b011111001111: data = 6'b010101;
12'b011111010000: data = 6'b010101;
12'b011111010001: data = 6'b010101;
12'b011111010010: data = 6'b010101;
12'b011111010011: data = 6'b010101;
12'b011111010100: data = 6'b010101;
12'b011111010101: data = 6'b010101;
12'b011111010110: data = 6'b010101;
12'b011111010111: data = 6'b010101;
12'b011111011000: data = 6'b010101;
12'b011111011001: data = 6'b101010;
12'b011111011010: data = 6'b101010;
12'b011111011011: data = 6'b101010;
12'b011111011100: data = 6'b101010;
12'b011111011101: data = 6'b101010;
12'b011111011110: data = 6'b101010;
12'b011111011111: data = 6'b101010;
12'b011111100000: data = 6'b010101;
12'b011111100001: data = 6'b010101;
12'b011111100010: data = 6'b010101;
12'b011111100011: data = 6'b010101;
12'b011111100100: data = 6'b010101;
12'b011111100101: data = 6'b010101;
12'b011111100110: data = 6'b010101;
12'b011111100111: data = 6'b000000;
12'b011111101000: data = 6'b000000;
12'b011111101001: data = 6'b000000;
12'b011111101010: data = 6'b000000;
12'b011111101011: data = 6'b000000;
12'b011111101100: data = 6'b000000;
12'b011111101101: data = 6'b000000;
12'b011111101110: data = 6'b000000;
12'b011111101111: data = 6'b000000;
12'b011111110000: data = 6'b000000;
12'b011111110001: data = 6'b000000;
12'b011111110010: data = 6'b000000;
12'b011111110011: data = 6'b000000;
12'b011111110100: data = 6'b000000;
12'b011111110101: data = 6'b000000;
12'b011111110110: data = 6'b000000;
12'b011111110111: data = 6'b000000;
12'b011111111000: data = 6'b000000;
12'b011111111001: data = 6'b000000;
12'b011111111010: data = 6'b000000;
12'b011111111011: data = 6'b000000;
12'b011111111100: data = 6'b000000;
12'b011111111101: data = 6'b000000;
12'b011111111110: data = 6'b000000;
12'b011111111111: data = 6'b000000;
12'b0111111000000: data = 6'b000000;
12'b0111111000001: data = 6'b000000;
12'b0111111000010: data = 6'b000000;
12'b0111111000011: data = 6'b000000;
12'b0111111000100: data = 6'b000000;
12'b0111111000101: data = 6'b000000;
12'b0111111000110: data = 6'b000000;
12'b0111111000111: data = 6'b000000;
12'b0111111001000: data = 6'b000000;
12'b0111111001001: data = 6'b000000;
12'b0111111001010: data = 6'b000000;
12'b0111111001011: data = 6'b000000;
12'b0111111001100: data = 6'b000000;
12'b0111111001101: data = 6'b000000;
12'b0111111001110: data = 6'b000000;
12'b0111111001111: data = 6'b000000;
12'b0111111010000: data = 6'b000000;
12'b0111111010001: data = 6'b000000;
12'b0111111010010: data = 6'b000000;
12'b0111111010011: data = 6'b000000;
12'b0111111010100: data = 6'b000000;
12'b0111111010101: data = 6'b000000;
12'b0111111010110: data = 6'b000000;
12'b0111111010111: data = 6'b000000;
12'b0111111011000: data = 6'b000000;
12'b0111111011001: data = 6'b000000;
12'b0111111011010: data = 6'b000000;
12'b0111111011011: data = 6'b000000;
12'b0111111011100: data = 6'b000000;
12'b0111111011101: data = 6'b000000;
12'b0111111011110: data = 6'b000000;
12'b0111111011111: data = 6'b000000;
12'b0111111100000: data = 6'b000000;
12'b0111111100001: data = 6'b000000;
12'b0111111100010: data = 6'b000000;
12'b0111111100011: data = 6'b000000;
12'b0111111100100: data = 6'b000000;
12'b0111111100101: data = 6'b000000;
12'b0111111100110: data = 6'b000000;
12'b0111111100111: data = 6'b000000;
12'b0111111101000: data = 6'b000000;
12'b0111111101001: data = 6'b000000;
12'b0111111101010: data = 6'b000000;
12'b0111111101011: data = 6'b000000;
12'b0111111101100: data = 6'b000000;
12'b0111111101101: data = 6'b000000;
12'b0111111101110: data = 6'b000000;
12'b0111111101111: data = 6'b000000;
12'b0111111110000: data = 6'b000000;
12'b0111111110001: data = 6'b000000;
12'b0111111110010: data = 6'b000000;
12'b0111111110011: data = 6'b000000;
12'b0111111110100: data = 6'b000000;
12'b0111111110101: data = 6'b000000;
12'b0111111110110: data = 6'b000000;
12'b0111111110111: data = 6'b000000;
12'b0111111111000: data = 6'b000000;
12'b0111111111001: data = 6'b000000;
12'b0111111111010: data = 6'b000000;
12'b0111111111011: data = 6'b000000;
12'b0111111111100: data = 6'b000000;
12'b0111111111101: data = 6'b000000;
12'b0111111111110: data = 6'b000000;
12'b0111111111111: data = 6'b000000;
12'b01111110000000: data = 6'b000000;
12'b01111110000001: data = 6'b000000;
12'b01111110000010: data = 6'b000000;
12'b01111110000011: data = 6'b000000;
12'b01111110000100: data = 6'b000000;
12'b01111110000101: data = 6'b000000;
12'b01111110000110: data = 6'b010101;
12'b01111110000111: data = 6'b010101;
12'b01111110001000: data = 6'b010101;
12'b01111110001001: data = 6'b010101;
12'b01111110001010: data = 6'b010101;
12'b01111110001011: data = 6'b101010;
12'b01111110001100: data = 6'b111111;
12'b01111110001101: data = 6'b101010;
12'b01111110001110: data = 6'b101010;
12'b01111110001111: data = 6'b101010;
12'b01111110010000: data = 6'b101010;
12'b01111110010001: data = 6'b101010;
12'b01111110010010: data = 6'b010101;
12'b01111110010011: data = 6'b010101;
12'b01111110010100: data = 6'b010101;
12'b01111110010101: data = 6'b010101;
12'b01111110010110: data = 6'b010101;
12'b01111110010111: data = 6'b010101;
12'b01111110011000: data = 6'b010101;
12'b01111110011001: data = 6'b010101;
12'b01111110011010: data = 6'b010101;
12'b01111110011011: data = 6'b010101;
12'b01111110011100: data = 6'b010101;
12'b01111110011101: data = 6'b010101;
12'b01111110011110: data = 6'b010101;
12'b01111110011111: data = 6'b010101;
12'b01111110100000: data = 6'b010101;
12'b01111110100001: data = 6'b010101;
12'b01111110100010: data = 6'b010101;
12'b01111110100011: data = 6'b010101;
12'b01111110100100: data = 6'b010101;
12'b01111110100101: data = 6'b010101;
12'b01111110100110: data = 6'b010101;
12'b01111110100111: data = 6'b010101;
12'b01111110101000: data = 6'b010101;
12'b01111110101001: data = 6'b010101;
12'b01111110101010: data = 6'b010101;
12'b100000000000: data = 6'b010101;
12'b100000000001: data = 6'b010101;
12'b100000000010: data = 6'b010101;
12'b100000000011: data = 6'b010101;
12'b100000000100: data = 6'b010101;
12'b100000000101: data = 6'b010101;
12'b100000000110: data = 6'b010101;
12'b100000000111: data = 6'b010101;
12'b100000001000: data = 6'b010101;
12'b100000001001: data = 6'b010101;
12'b100000001010: data = 6'b010101;
12'b100000001011: data = 6'b010101;
12'b100000001100: data = 6'b010101;
12'b100000001101: data = 6'b010101;
12'b100000001110: data = 6'b010101;
12'b100000001111: data = 6'b010101;
12'b100000010000: data = 6'b010101;
12'b100000010001: data = 6'b010101;
12'b100000010010: data = 6'b010101;
12'b100000010011: data = 6'b010101;
12'b100000010100: data = 6'b010101;
12'b100000010101: data = 6'b010101;
12'b100000010110: data = 6'b010101;
12'b100000010111: data = 6'b010101;
12'b100000011000: data = 6'b010101;
12'b100000011001: data = 6'b101010;
12'b100000011010: data = 6'b101010;
12'b100000011011: data = 6'b101010;
12'b100000011100: data = 6'b101010;
12'b100000011101: data = 6'b101010;
12'b100000011110: data = 6'b101010;
12'b100000011111: data = 6'b101010;
12'b100000100000: data = 6'b010101;
12'b100000100001: data = 6'b010101;
12'b100000100010: data = 6'b010101;
12'b100000100011: data = 6'b010101;
12'b100000100100: data = 6'b010101;
12'b100000100101: data = 6'b010101;
12'b100000100110: data = 6'b010101;
12'b100000100111: data = 6'b000000;
12'b100000101000: data = 6'b000000;
12'b100000101001: data = 6'b000000;
12'b100000101010: data = 6'b000000;
12'b100000101011: data = 6'b000000;
12'b100000101100: data = 6'b000000;
12'b100000101101: data = 6'b000000;
12'b100000101110: data = 6'b000000;
12'b100000101111: data = 6'b000000;
12'b100000110000: data = 6'b000000;
12'b100000110001: data = 6'b000000;
12'b100000110010: data = 6'b000000;
12'b100000110011: data = 6'b000000;
12'b100000110100: data = 6'b000000;
12'b100000110101: data = 6'b000000;
12'b100000110110: data = 6'b000000;
12'b100000110111: data = 6'b000000;
12'b100000111000: data = 6'b000000;
12'b100000111001: data = 6'b000000;
12'b100000111010: data = 6'b000000;
12'b100000111011: data = 6'b000000;
12'b100000111100: data = 6'b000000;
12'b100000111101: data = 6'b000000;
12'b100000111110: data = 6'b000000;
12'b100000111111: data = 6'b000000;
12'b1000001000000: data = 6'b000000;
12'b1000001000001: data = 6'b000000;
12'b1000001000010: data = 6'b000000;
12'b1000001000011: data = 6'b000000;
12'b1000001000100: data = 6'b000000;
12'b1000001000101: data = 6'b000000;
12'b1000001000110: data = 6'b000000;
12'b1000001000111: data = 6'b000000;
12'b1000001001000: data = 6'b000000;
12'b1000001001001: data = 6'b000000;
12'b1000001001010: data = 6'b000000;
12'b1000001001011: data = 6'b000000;
12'b1000001001100: data = 6'b000000;
12'b1000001001101: data = 6'b000000;
12'b1000001001110: data = 6'b000000;
12'b1000001001111: data = 6'b000000;
12'b1000001010000: data = 6'b000000;
12'b1000001010001: data = 6'b000000;
12'b1000001010010: data = 6'b000000;
12'b1000001010011: data = 6'b000000;
12'b1000001010100: data = 6'b000000;
12'b1000001010101: data = 6'b000000;
12'b1000001010110: data = 6'b000000;
12'b1000001010111: data = 6'b000000;
12'b1000001011000: data = 6'b000000;
12'b1000001011001: data = 6'b000000;
12'b1000001011010: data = 6'b000000;
12'b1000001011011: data = 6'b000000;
12'b1000001011100: data = 6'b000000;
12'b1000001011101: data = 6'b000000;
12'b1000001011110: data = 6'b000000;
12'b1000001011111: data = 6'b000000;
12'b1000001100000: data = 6'b000000;
12'b1000001100001: data = 6'b000000;
12'b1000001100010: data = 6'b000000;
12'b1000001100011: data = 6'b000000;
12'b1000001100100: data = 6'b000000;
12'b1000001100101: data = 6'b000000;
12'b1000001100110: data = 6'b000000;
12'b1000001100111: data = 6'b000000;
12'b1000001101000: data = 6'b000000;
12'b1000001101001: data = 6'b000000;
12'b1000001101010: data = 6'b000000;
12'b1000001101011: data = 6'b000000;
12'b1000001101100: data = 6'b000000;
12'b1000001101101: data = 6'b000000;
12'b1000001101110: data = 6'b000000;
12'b1000001101111: data = 6'b000000;
12'b1000001110000: data = 6'b000000;
12'b1000001110001: data = 6'b000000;
12'b1000001110010: data = 6'b000000;
12'b1000001110011: data = 6'b000000;
12'b1000001110100: data = 6'b000000;
12'b1000001110101: data = 6'b000000;
12'b1000001110110: data = 6'b000000;
12'b1000001110111: data = 6'b000000;
12'b1000001111000: data = 6'b000000;
12'b1000001111001: data = 6'b000000;
12'b1000001111010: data = 6'b000000;
12'b1000001111011: data = 6'b000000;
12'b1000001111100: data = 6'b000000;
12'b1000001111101: data = 6'b000000;
12'b1000001111110: data = 6'b000000;
12'b1000001111111: data = 6'b000000;
12'b10000010000000: data = 6'b000000;
12'b10000010000001: data = 6'b000000;
12'b10000010000010: data = 6'b000000;
12'b10000010000011: data = 6'b000000;
12'b10000010000100: data = 6'b000000;
12'b10000010000101: data = 6'b010101;
12'b10000010000110: data = 6'b010101;
12'b10000010000111: data = 6'b010101;
12'b10000010001000: data = 6'b010101;
12'b10000010001001: data = 6'b010101;
12'b10000010001010: data = 6'b010101;
12'b10000010001011: data = 6'b101010;
12'b10000010001100: data = 6'b101010;
12'b10000010001101: data = 6'b101010;
12'b10000010001110: data = 6'b101010;
12'b10000010001111: data = 6'b101010;
12'b10000010010000: data = 6'b101010;
12'b10000010010001: data = 6'b101010;
12'b10000010010010: data = 6'b010101;
12'b10000010010011: data = 6'b010101;
12'b10000010010100: data = 6'b010101;
12'b10000010010101: data = 6'b010101;
12'b10000010010110: data = 6'b010101;
12'b10000010010111: data = 6'b010101;
12'b10000010011000: data = 6'b010101;
12'b10000010011001: data = 6'b010101;
12'b10000010011010: data = 6'b010101;
12'b10000010011011: data = 6'b010101;
12'b10000010011100: data = 6'b010101;
12'b10000010011101: data = 6'b010101;
12'b10000010011110: data = 6'b010101;
12'b10000010011111: data = 6'b010101;
12'b10000010100000: data = 6'b010101;
12'b10000010100001: data = 6'b010101;
12'b10000010100010: data = 6'b010101;
12'b10000010100011: data = 6'b010101;
12'b10000010100100: data = 6'b010101;
12'b10000010100101: data = 6'b010101;
12'b10000010100110: data = 6'b010101;
12'b10000010100111: data = 6'b010101;
12'b10000010101000: data = 6'b010101;
12'b10000010101001: data = 6'b010101;
12'b10000010101010: data = 6'b010101;
12'b100001000000: data = 6'b010101;
12'b100001000001: data = 6'b010101;
12'b100001000010: data = 6'b010101;
12'b100001000011: data = 6'b010101;
12'b100001000100: data = 6'b010101;
12'b100001000101: data = 6'b010101;
12'b100001000110: data = 6'b010101;
12'b100001000111: data = 6'b010101;
12'b100001001000: data = 6'b010101;
12'b100001001001: data = 6'b010101;
12'b100001001010: data = 6'b010101;
12'b100001001011: data = 6'b010101;
12'b100001001100: data = 6'b010101;
12'b100001001101: data = 6'b010101;
12'b100001001110: data = 6'b010101;
12'b100001001111: data = 6'b010101;
12'b100001010000: data = 6'b010101;
12'b100001010001: data = 6'b010101;
12'b100001010010: data = 6'b010101;
12'b100001010011: data = 6'b010101;
12'b100001010100: data = 6'b010101;
12'b100001010101: data = 6'b010101;
12'b100001010110: data = 6'b010101;
12'b100001010111: data = 6'b010101;
12'b100001011000: data = 6'b010101;
12'b100001011001: data = 6'b101010;
12'b100001011010: data = 6'b101010;
12'b100001011011: data = 6'b101010;
12'b100001011100: data = 6'b101010;
12'b100001011101: data = 6'b101010;
12'b100001011110: data = 6'b101010;
12'b100001011111: data = 6'b101010;
12'b100001100000: data = 6'b010101;
12'b100001100001: data = 6'b010101;
12'b100001100010: data = 6'b010101;
12'b100001100011: data = 6'b010101;
12'b100001100100: data = 6'b010101;
12'b100001100101: data = 6'b010101;
12'b100001100110: data = 6'b010101;
12'b100001100111: data = 6'b000000;
12'b100001101000: data = 6'b000000;
12'b100001101001: data = 6'b000000;
12'b100001101010: data = 6'b000000;
12'b100001101011: data = 6'b000000;
12'b100001101100: data = 6'b000000;
12'b100001101101: data = 6'b000000;
12'b100001101110: data = 6'b000000;
12'b100001101111: data = 6'b000000;
12'b100001110000: data = 6'b000000;
12'b100001110001: data = 6'b000000;
12'b100001110010: data = 6'b000000;
12'b100001110011: data = 6'b000000;
12'b100001110100: data = 6'b000000;
12'b100001110101: data = 6'b000000;
12'b100001110110: data = 6'b000000;
12'b100001110111: data = 6'b000000;
12'b100001111000: data = 6'b000000;
12'b100001111001: data = 6'b000000;
12'b100001111010: data = 6'b000000;
12'b100001111011: data = 6'b000000;
12'b100001111100: data = 6'b000000;
12'b100001111101: data = 6'b000000;
12'b100001111110: data = 6'b000000;
12'b100001111111: data = 6'b000000;
12'b1000011000000: data = 6'b000000;
12'b1000011000001: data = 6'b000000;
12'b1000011000010: data = 6'b000000;
12'b1000011000011: data = 6'b000000;
12'b1000011000100: data = 6'b000000;
12'b1000011000101: data = 6'b000000;
12'b1000011000110: data = 6'b000000;
12'b1000011000111: data = 6'b000000;
12'b1000011001000: data = 6'b000000;
12'b1000011001001: data = 6'b000000;
12'b1000011001010: data = 6'b000000;
12'b1000011001011: data = 6'b000000;
12'b1000011001100: data = 6'b000000;
12'b1000011001101: data = 6'b000000;
12'b1000011001110: data = 6'b000000;
12'b1000011001111: data = 6'b000000;
12'b1000011010000: data = 6'b000000;
12'b1000011010001: data = 6'b000000;
12'b1000011010010: data = 6'b000000;
12'b1000011010011: data = 6'b000000;
12'b1000011010100: data = 6'b000000;
12'b1000011010101: data = 6'b000000;
12'b1000011010110: data = 6'b000000;
12'b1000011010111: data = 6'b000000;
12'b1000011011000: data = 6'b000000;
12'b1000011011001: data = 6'b000000;
12'b1000011011010: data = 6'b000000;
12'b1000011011011: data = 6'b000000;
12'b1000011011100: data = 6'b000000;
12'b1000011011101: data = 6'b000000;
12'b1000011011110: data = 6'b000000;
12'b1000011011111: data = 6'b000000;
12'b1000011100000: data = 6'b000000;
12'b1000011100001: data = 6'b000000;
12'b1000011100010: data = 6'b000000;
12'b1000011100011: data = 6'b000000;
12'b1000011100100: data = 6'b000000;
12'b1000011100101: data = 6'b000000;
12'b1000011100110: data = 6'b000000;
12'b1000011100111: data = 6'b000000;
12'b1000011101000: data = 6'b000000;
12'b1000011101001: data = 6'b000000;
12'b1000011101010: data = 6'b000000;
12'b1000011101011: data = 6'b000000;
12'b1000011101100: data = 6'b000000;
12'b1000011101101: data = 6'b000000;
12'b1000011101110: data = 6'b000000;
12'b1000011101111: data = 6'b000000;
12'b1000011110000: data = 6'b000000;
12'b1000011110001: data = 6'b000000;
12'b1000011110010: data = 6'b000000;
12'b1000011110011: data = 6'b000000;
12'b1000011110100: data = 6'b000000;
12'b1000011110101: data = 6'b000000;
12'b1000011110110: data = 6'b000000;
12'b1000011110111: data = 6'b000000;
12'b1000011111000: data = 6'b000000;
12'b1000011111001: data = 6'b000000;
12'b1000011111010: data = 6'b000000;
12'b1000011111011: data = 6'b000000;
12'b1000011111100: data = 6'b000000;
12'b1000011111101: data = 6'b000000;
12'b1000011111110: data = 6'b000000;
12'b1000011111111: data = 6'b000000;
12'b10000110000000: data = 6'b000000;
12'b10000110000001: data = 6'b000000;
12'b10000110000010: data = 6'b000000;
12'b10000110000011: data = 6'b000000;
12'b10000110000100: data = 6'b000000;
12'b10000110000101: data = 6'b000000;
12'b10000110000110: data = 6'b010101;
12'b10000110000111: data = 6'b010101;
12'b10000110001000: data = 6'b010101;
12'b10000110001001: data = 6'b010101;
12'b10000110001010: data = 6'b010101;
12'b10000110001011: data = 6'b101010;
12'b10000110001100: data = 6'b101010;
12'b10000110001101: data = 6'b101010;
12'b10000110001110: data = 6'b101010;
12'b10000110001111: data = 6'b101010;
12'b10000110010000: data = 6'b101010;
12'b10000110010001: data = 6'b101010;
12'b10000110010010: data = 6'b010101;
12'b10000110010011: data = 6'b010101;
12'b10000110010100: data = 6'b010101;
12'b10000110010101: data = 6'b010101;
12'b10000110010110: data = 6'b010101;
12'b10000110010111: data = 6'b010101;
12'b10000110011000: data = 6'b010101;
12'b10000110011001: data = 6'b010101;
12'b10000110011010: data = 6'b010101;
12'b10000110011011: data = 6'b010101;
12'b10000110011100: data = 6'b010101;
12'b10000110011101: data = 6'b010101;
12'b10000110011110: data = 6'b010101;
12'b10000110011111: data = 6'b010101;
12'b10000110100000: data = 6'b010101;
12'b10000110100001: data = 6'b010101;
12'b10000110100010: data = 6'b010101;
12'b10000110100011: data = 6'b010101;
12'b10000110100100: data = 6'b010101;
12'b10000110100101: data = 6'b010101;
12'b10000110100110: data = 6'b010101;
12'b10000110100111: data = 6'b010101;
12'b10000110101000: data = 6'b010101;
12'b10000110101001: data = 6'b010101;
12'b10000110101010: data = 6'b010101;
12'b100010000000: data = 6'b010101;
12'b100010000001: data = 6'b010101;
12'b100010000010: data = 6'b010101;
12'b100010000011: data = 6'b010101;
12'b100010000100: data = 6'b010101;
12'b100010000101: data = 6'b010101;
12'b100010000110: data = 6'b010101;
12'b100010000111: data = 6'b010101;
12'b100010001000: data = 6'b010101;
12'b100010001001: data = 6'b010101;
12'b100010001010: data = 6'b010101;
12'b100010001011: data = 6'b010101;
12'b100010001100: data = 6'b010101;
12'b100010001101: data = 6'b010101;
12'b100010001110: data = 6'b010101;
12'b100010001111: data = 6'b010101;
12'b100010010000: data = 6'b010101;
12'b100010010001: data = 6'b010101;
12'b100010010010: data = 6'b010101;
12'b100010010011: data = 6'b010101;
12'b100010010100: data = 6'b010101;
12'b100010010101: data = 6'b010101;
12'b100010010110: data = 6'b010101;
12'b100010010111: data = 6'b010101;
12'b100010011000: data = 6'b010101;
12'b100010011001: data = 6'b101010;
12'b100010011010: data = 6'b101010;
12'b100010011011: data = 6'b101010;
12'b100010011100: data = 6'b101010;
12'b100010011101: data = 6'b010101;
12'b100010011110: data = 6'b010101;
12'b100010011111: data = 6'b010101;
12'b100010100000: data = 6'b010101;
12'b100010100001: data = 6'b010101;
12'b100010100010: data = 6'b010101;
12'b100010100011: data = 6'b010101;
12'b100010100100: data = 6'b010101;
12'b100010100101: data = 6'b010101;
12'b100010100110: data = 6'b010101;
12'b100010100111: data = 6'b010101;
12'b100010101000: data = 6'b010101;
12'b100010101001: data = 6'b010101;
12'b100010101010: data = 6'b010101;
12'b100010101011: data = 6'b010101;
12'b100010101100: data = 6'b010101;
12'b100010101101: data = 6'b010101;
12'b100010101110: data = 6'b010101;
12'b100010101111: data = 6'b010101;
12'b100010110000: data = 6'b010101;
12'b100010110001: data = 6'b010101;
12'b100010110010: data = 6'b010101;
12'b100010110011: data = 6'b010101;
12'b100010110100: data = 6'b010101;
12'b100010110101: data = 6'b010101;
12'b100010110110: data = 6'b010101;
12'b100010110111: data = 6'b010101;
12'b100010111000: data = 6'b010101;
12'b100010111001: data = 6'b010101;
12'b100010111010: data = 6'b010101;
12'b100010111011: data = 6'b010101;
12'b100010111100: data = 6'b010101;
12'b100010111101: data = 6'b010101;
12'b100010111110: data = 6'b010101;
12'b100010111111: data = 6'b010101;
12'b1000101000000: data = 6'b010101;
12'b1000101000001: data = 6'b010101;
12'b1000101000010: data = 6'b010101;
12'b1000101000011: data = 6'b010101;
12'b1000101000100: data = 6'b010101;
12'b1000101000101: data = 6'b010101;
12'b1000101000110: data = 6'b010101;
12'b1000101000111: data = 6'b010101;
12'b1000101001000: data = 6'b010101;
12'b1000101001001: data = 6'b010101;
12'b1000101001010: data = 6'b010101;
12'b1000101001011: data = 6'b010101;
12'b1000101001100: data = 6'b010101;
12'b1000101001101: data = 6'b010101;
12'b1000101001110: data = 6'b010101;
12'b1000101001111: data = 6'b010101;
12'b1000101010000: data = 6'b010101;
12'b1000101010001: data = 6'b010101;
12'b1000101010010: data = 6'b010101;
12'b1000101010011: data = 6'b010101;
12'b1000101010100: data = 6'b010101;
12'b1000101010101: data = 6'b010101;
12'b1000101010110: data = 6'b010101;
12'b1000101010111: data = 6'b010101;
12'b1000101011000: data = 6'b010101;
12'b1000101011001: data = 6'b010101;
12'b1000101011010: data = 6'b010101;
12'b1000101011011: data = 6'b010101;
12'b1000101011100: data = 6'b010101;
12'b1000101011101: data = 6'b010101;
12'b1000101011110: data = 6'b010101;
12'b1000101011111: data = 6'b010101;
12'b1000101100000: data = 6'b010101;
12'b1000101100001: data = 6'b010101;
12'b1000101100010: data = 6'b010101;
12'b1000101100011: data = 6'b010101;
12'b1000101100100: data = 6'b010101;
12'b1000101100101: data = 6'b010101;
12'b1000101100110: data = 6'b010101;
12'b1000101100111: data = 6'b010101;
12'b1000101101000: data = 6'b010101;
12'b1000101101001: data = 6'b010101;
12'b1000101101010: data = 6'b010101;
12'b1000101101011: data = 6'b010101;
12'b1000101101100: data = 6'b010101;
12'b1000101101101: data = 6'b010101;
12'b1000101101110: data = 6'b010101;
12'b1000101101111: data = 6'b010101;
12'b1000101110000: data = 6'b010101;
12'b1000101110001: data = 6'b010101;
12'b1000101110010: data = 6'b010101;
12'b1000101110011: data = 6'b010101;
12'b1000101110100: data = 6'b010101;
12'b1000101110101: data = 6'b010101;
12'b1000101110110: data = 6'b010101;
12'b1000101110111: data = 6'b010101;
12'b1000101111000: data = 6'b010101;
12'b1000101111001: data = 6'b010101;
12'b1000101111010: data = 6'b010101;
12'b1000101111011: data = 6'b010101;
12'b1000101111100: data = 6'b010101;
12'b1000101111101: data = 6'b010101;
12'b1000101111110: data = 6'b010101;
12'b1000101111111: data = 6'b010101;
12'b10001010000000: data = 6'b010101;
12'b10001010000001: data = 6'b010101;
12'b10001010000010: data = 6'b010101;
12'b10001010000011: data = 6'b010101;
12'b10001010000100: data = 6'b010101;
12'b10001010000101: data = 6'b010101;
12'b10001010000110: data = 6'b010101;
12'b10001010000111: data = 6'b010101;
12'b10001010001000: data = 6'b010101;
12'b10001010001001: data = 6'b010101;
12'b10001010001010: data = 6'b010101;
12'b10001010001011: data = 6'b010101;
12'b10001010001100: data = 6'b101001;
12'b10001010001101: data = 6'b101001;
12'b10001010001110: data = 6'b101010;
12'b10001010001111: data = 6'b101010;
12'b10001010010000: data = 6'b101010;
12'b10001010010001: data = 6'b101010;
12'b10001010010010: data = 6'b010101;
12'b10001010010011: data = 6'b010101;
12'b10001010010100: data = 6'b010101;
12'b10001010010101: data = 6'b010101;
12'b10001010010110: data = 6'b010101;
12'b10001010010111: data = 6'b010101;
12'b10001010011000: data = 6'b010101;
12'b10001010011001: data = 6'b010101;
12'b10001010011010: data = 6'b010101;
12'b10001010011011: data = 6'b010101;
12'b10001010011100: data = 6'b010101;
12'b10001010011101: data = 6'b010101;
12'b10001010011110: data = 6'b010101;
12'b10001010011111: data = 6'b010101;
12'b10001010100000: data = 6'b010101;
12'b10001010100001: data = 6'b010101;
12'b10001010100010: data = 6'b010101;
12'b10001010100011: data = 6'b010101;
12'b10001010100100: data = 6'b010101;
12'b10001010100101: data = 6'b010101;
12'b10001010100110: data = 6'b010101;
12'b10001010100111: data = 6'b010101;
12'b10001010101000: data = 6'b010101;
12'b10001010101001: data = 6'b010101;
12'b10001010101010: data = 6'b010101;
12'b100011000000: data = 6'b010101;
12'b100011000001: data = 6'b010101;
12'b100011000010: data = 6'b010101;
12'b100011000011: data = 6'b010101;
12'b100011000100: data = 6'b010101;
12'b100011000101: data = 6'b010101;
12'b100011000110: data = 6'b010101;
12'b100011000111: data = 6'b010101;
12'b100011001000: data = 6'b010101;
12'b100011001001: data = 6'b010101;
12'b100011001010: data = 6'b010101;
12'b100011001011: data = 6'b010101;
12'b100011001100: data = 6'b010101;
12'b100011001101: data = 6'b010101;
12'b100011001110: data = 6'b010101;
12'b100011001111: data = 6'b010101;
12'b100011010000: data = 6'b010101;
12'b100011010001: data = 6'b010101;
12'b100011010010: data = 6'b010101;
12'b100011010011: data = 6'b010101;
12'b100011010100: data = 6'b010101;
12'b100011010101: data = 6'b010101;
12'b100011010110: data = 6'b010101;
12'b100011010111: data = 6'b010101;
12'b100011011000: data = 6'b010101;
12'b100011011001: data = 6'b101010;
12'b100011011010: data = 6'b101010;
12'b100011011011: data = 6'b101010;
12'b100011011100: data = 6'b010101;
12'b100011011101: data = 6'b000000;
12'b100011011110: data = 6'b000000;
12'b100011011111: data = 6'b010101;
12'b100011100000: data = 6'b010101;
12'b100011100001: data = 6'b010101;
12'b100011100010: data = 6'b010101;
12'b100011100011: data = 6'b010101;
12'b100011100100: data = 6'b010101;
12'b100011100101: data = 6'b101001;
12'b100011100110: data = 6'b101010;
12'b100011100111: data = 6'b101010;
12'b100011101000: data = 6'b101010;
12'b100011101001: data = 6'b101010;
12'b100011101010: data = 6'b101010;
12'b100011101011: data = 6'b101010;
12'b100011101100: data = 6'b101010;
12'b100011101101: data = 6'b101010;
12'b100011101110: data = 6'b101010;
12'b100011101111: data = 6'b101010;
12'b100011110000: data = 6'b101010;
12'b100011110001: data = 6'b101010;
12'b100011110010: data = 6'b101010;
12'b100011110011: data = 6'b101010;
12'b100011110100: data = 6'b101010;
12'b100011110101: data = 6'b111010;
12'b100011110110: data = 6'b111010;
12'b100011110111: data = 6'b111110;
12'b100011111000: data = 6'b111111;
12'b100011111001: data = 6'b111111;
12'b100011111010: data = 6'b111111;
12'b100011111011: data = 6'b111111;
12'b100011111100: data = 6'b111111;
12'b100011111101: data = 6'b111111;
12'b100011111110: data = 6'b111111;
12'b100011111111: data = 6'b111111;
12'b1000111000000: data = 6'b111111;
12'b1000111000001: data = 6'b111111;
12'b1000111000010: data = 6'b111111;
12'b1000111000011: data = 6'b111111;
12'b1000111000100: data = 6'b111111;
12'b1000111000101: data = 6'b111111;
12'b1000111000110: data = 6'b111111;
12'b1000111000111: data = 6'b111110;
12'b1000111001000: data = 6'b111110;
12'b1000111001001: data = 6'b111110;
12'b1000111001010: data = 6'b111110;
12'b1000111001011: data = 6'b111110;
12'b1000111001100: data = 6'b111010;
12'b1000111001101: data = 6'b111010;
12'b1000111001110: data = 6'b111010;
12'b1000111001111: data = 6'b101010;
12'b1000111010000: data = 6'b101010;
12'b1000111010001: data = 6'b101010;
12'b1000111010010: data = 6'b101010;
12'b1000111010011: data = 6'b101010;
12'b1000111010100: data = 6'b101010;
12'b1000111010101: data = 6'b101010;
12'b1000111010110: data = 6'b101010;
12'b1000111010111: data = 6'b101010;
12'b1000111011000: data = 6'b101010;
12'b1000111011001: data = 6'b101010;
12'b1000111011010: data = 6'b101010;
12'b1000111011011: data = 6'b101010;
12'b1000111011100: data = 6'b101010;
12'b1000111011101: data = 6'b101010;
12'b1000111011110: data = 6'b101010;
12'b1000111011111: data = 6'b101010;
12'b1000111100000: data = 6'b101010;
12'b1000111100001: data = 6'b101010;
12'b1000111100010: data = 6'b101010;
12'b1000111100011: data = 6'b101010;
12'b1000111100100: data = 6'b101010;
12'b1000111100101: data = 6'b101010;
12'b1000111100110: data = 6'b101010;
12'b1000111100111: data = 6'b101010;
12'b1000111101000: data = 6'b101010;
12'b1000111101001: data = 6'b101010;
12'b1000111101010: data = 6'b101010;
12'b1000111101011: data = 6'b101010;
12'b1000111101100: data = 6'b101010;
12'b1000111101101: data = 6'b101010;
12'b1000111101110: data = 6'b101010;
12'b1000111101111: data = 6'b101010;
12'b1000111110000: data = 6'b101010;
12'b1000111110001: data = 6'b101010;
12'b1000111110010: data = 6'b101010;
12'b1000111110011: data = 6'b101010;
12'b1000111110100: data = 6'b101010;
12'b1000111110101: data = 6'b101010;
12'b1000111110110: data = 6'b101010;
12'b1000111110111: data = 6'b101010;
12'b1000111111000: data = 6'b101010;
12'b1000111111001: data = 6'b101010;
12'b1000111111010: data = 6'b101010;
12'b1000111111011: data = 6'b101001;
12'b1000111111100: data = 6'b101001;
12'b1000111111101: data = 6'b101001;
12'b1000111111110: data = 6'b101001;
12'b1000111111111: data = 6'b010101;
12'b10001110000000: data = 6'b010101;
12'b10001110000001: data = 6'b010101;
12'b10001110000010: data = 6'b010101;
12'b10001110000011: data = 6'b010101;
12'b10001110000100: data = 6'b010101;
12'b10001110000101: data = 6'b010101;
12'b10001110000110: data = 6'b010101;
12'b10001110000111: data = 6'b010101;
12'b10001110001000: data = 6'b010101;
12'b10001110001001: data = 6'b010101;
12'b10001110001010: data = 6'b010101;
12'b10001110001011: data = 6'b010101;
12'b10001110001100: data = 6'b000000;
12'b10001110001101: data = 6'b000000;
12'b10001110001110: data = 6'b101010;
12'b10001110001111: data = 6'b101010;
12'b10001110010000: data = 6'b101010;
12'b10001110010001: data = 6'b101010;
12'b10001110010010: data = 6'b010101;
12'b10001110010011: data = 6'b010101;
12'b10001110010100: data = 6'b010101;
12'b10001110010101: data = 6'b010101;
12'b10001110010110: data = 6'b010101;
12'b10001110010111: data = 6'b010101;
12'b10001110011000: data = 6'b010101;
12'b10001110011001: data = 6'b010101;
12'b10001110011010: data = 6'b010101;
12'b10001110011011: data = 6'b010101;
12'b10001110011100: data = 6'b010101;
12'b10001110011101: data = 6'b010101;
12'b10001110011110: data = 6'b010101;
12'b10001110011111: data = 6'b010101;
12'b10001110100000: data = 6'b010101;
12'b10001110100001: data = 6'b010101;
12'b10001110100010: data = 6'b010101;
12'b10001110100011: data = 6'b010101;
12'b10001110100100: data = 6'b010101;
12'b10001110100101: data = 6'b010101;
12'b10001110100110: data = 6'b010101;
12'b10001110100111: data = 6'b010101;
12'b10001110101000: data = 6'b010101;
12'b10001110101001: data = 6'b010101;
12'b10001110101010: data = 6'b010101;
12'b100100000000: data = 6'b010101;
12'b100100000001: data = 6'b010101;
12'b100100000010: data = 6'b010101;
12'b100100000011: data = 6'b010101;
12'b100100000100: data = 6'b010101;
12'b100100000101: data = 6'b010101;
12'b100100000110: data = 6'b010101;
12'b100100000111: data = 6'b010101;
12'b100100001000: data = 6'b010101;
12'b100100001001: data = 6'b010101;
12'b100100001010: data = 6'b010101;
12'b100100001011: data = 6'b010101;
12'b100100001100: data = 6'b010101;
12'b100100001101: data = 6'b010101;
12'b100100001110: data = 6'b010101;
12'b100100001111: data = 6'b010101;
12'b100100010000: data = 6'b010101;
12'b100100010001: data = 6'b010101;
12'b100100010010: data = 6'b010101;
12'b100100010011: data = 6'b010101;
12'b100100010100: data = 6'b010101;
12'b100100010101: data = 6'b010101;
12'b100100010110: data = 6'b010101;
12'b100100010111: data = 6'b010101;
12'b100100011000: data = 6'b010101;
12'b100100011001: data = 6'b101010;
12'b100100011010: data = 6'b101010;
12'b100100011011: data = 6'b101010;
12'b100100011100: data = 6'b010101;
12'b100100011101: data = 6'b000000;
12'b100100011110: data = 6'b000000;
12'b100100011111: data = 6'b010101;
12'b100100100000: data = 6'b010101;
12'b100100100001: data = 6'b010101;
12'b100100100010: data = 6'b010101;
12'b100100100011: data = 6'b010101;
12'b100100100100: data = 6'b010101;
12'b100100100101: data = 6'b101001;
12'b100100100110: data = 6'b101001;
12'b100100100111: data = 6'b101010;
12'b100100101000: data = 6'b101010;
12'b100100101001: data = 6'b101010;
12'b100100101010: data = 6'b101010;
12'b100100101011: data = 6'b101010;
12'b100100101100: data = 6'b101010;
12'b100100101101: data = 6'b101010;
12'b100100101110: data = 6'b101010;
12'b100100101111: data = 6'b101010;
12'b100100110000: data = 6'b101010;
12'b100100110001: data = 6'b101010;
12'b100100110010: data = 6'b101010;
12'b100100110011: data = 6'b101010;
12'b100100110100: data = 6'b101010;
12'b100100110101: data = 6'b111010;
12'b100100110110: data = 6'b111010;
12'b100100110111: data = 6'b111110;
12'b100100111000: data = 6'b111110;
12'b100100111001: data = 6'b111111;
12'b100100111010: data = 6'b111111;
12'b100100111011: data = 6'b111111;
12'b100100111100: data = 6'b111111;
12'b100100111101: data = 6'b111111;
12'b100100111110: data = 6'b111111;
12'b100100111111: data = 6'b111111;
12'b1001001000000: data = 6'b111111;
12'b1001001000001: data = 6'b111111;
12'b1001001000010: data = 6'b111111;
12'b1001001000011: data = 6'b111111;
12'b1001001000100: data = 6'b111111;
12'b1001001000101: data = 6'b111111;
12'b1001001000110: data = 6'b111111;
12'b1001001000111: data = 6'b111110;
12'b1001001001000: data = 6'b111110;
12'b1001001001001: data = 6'b111110;
12'b1001001001010: data = 6'b111110;
12'b1001001001011: data = 6'b111110;
12'b1001001001100: data = 6'b111010;
12'b1001001001101: data = 6'b111010;
12'b1001001001110: data = 6'b111010;
12'b1001001001111: data = 6'b101010;
12'b1001001010000: data = 6'b101010;
12'b1001001010001: data = 6'b101010;
12'b1001001010010: data = 6'b101010;
12'b1001001010011: data = 6'b101010;
12'b1001001010100: data = 6'b101010;
12'b1001001010101: data = 6'b101010;
12'b1001001010110: data = 6'b101010;
12'b1001001010111: data = 6'b101010;
12'b1001001011000: data = 6'b101010;
12'b1001001011001: data = 6'b101010;
12'b1001001011010: data = 6'b101010;
12'b1001001011011: data = 6'b101010;
12'b1001001011100: data = 6'b101010;
12'b1001001011101: data = 6'b101010;
12'b1001001011110: data = 6'b101010;
12'b1001001011111: data = 6'b101010;
12'b1001001100000: data = 6'b101010;
12'b1001001100001: data = 6'b101010;
12'b1001001100010: data = 6'b101010;
12'b1001001100011: data = 6'b101010;
12'b1001001100100: data = 6'b101010;
12'b1001001100101: data = 6'b101010;
12'b1001001100110: data = 6'b101010;
12'b1001001100111: data = 6'b101010;
12'b1001001101000: data = 6'b101010;
12'b1001001101001: data = 6'b101010;
12'b1001001101010: data = 6'b101010;
12'b1001001101011: data = 6'b101010;
12'b1001001101100: data = 6'b101010;
12'b1001001101101: data = 6'b101010;
12'b1001001101110: data = 6'b101010;
12'b1001001101111: data = 6'b101010;
12'b1001001110000: data = 6'b101010;
12'b1001001110001: data = 6'b101010;
12'b1001001110010: data = 6'b101010;
12'b1001001110011: data = 6'b101010;
12'b1001001110100: data = 6'b101010;
12'b1001001110101: data = 6'b101010;
12'b1001001110110: data = 6'b101010;
12'b1001001110111: data = 6'b101010;
12'b1001001111000: data = 6'b101010;
12'b1001001111001: data = 6'b101001;
12'b1001001111010: data = 6'b101001;
12'b1001001111011: data = 6'b101001;
12'b1001001111100: data = 6'b101001;
12'b1001001111101: data = 6'b101001;
12'b1001001111110: data = 6'b010101;
12'b1001001111111: data = 6'b010101;
12'b10010010000000: data = 6'b010101;
12'b10010010000001: data = 6'b010101;
12'b10010010000010: data = 6'b010101;
12'b10010010000011: data = 6'b010101;
12'b10010010000100: data = 6'b010101;
12'b10010010000101: data = 6'b010101;
12'b10010010000110: data = 6'b010101;
12'b10010010000111: data = 6'b010101;
12'b10010010001000: data = 6'b010101;
12'b10010010001001: data = 6'b010101;
12'b10010010001010: data = 6'b010101;
12'b10010010001011: data = 6'b010101;
12'b10010010001100: data = 6'b000000;
12'b10010010001101: data = 6'b000000;
12'b10010010001110: data = 6'b101010;
12'b10010010001111: data = 6'b101010;
12'b10010010010000: data = 6'b101010;
12'b10010010010001: data = 6'b101010;
12'b10010010010010: data = 6'b010101;
12'b10010010010011: data = 6'b010101;
12'b10010010010100: data = 6'b010101;
12'b10010010010101: data = 6'b010101;
12'b10010010010110: data = 6'b010101;
12'b10010010010111: data = 6'b010101;
12'b10010010011000: data = 6'b010101;
12'b10010010011001: data = 6'b010101;
12'b10010010011010: data = 6'b010101;
12'b10010010011011: data = 6'b010101;
12'b10010010011100: data = 6'b010101;
12'b10010010011101: data = 6'b010101;
12'b10010010011110: data = 6'b010101;
12'b10010010011111: data = 6'b010101;
12'b10010010100000: data = 6'b010101;
12'b10010010100001: data = 6'b010101;
12'b10010010100010: data = 6'b010101;
12'b10010010100011: data = 6'b010101;
12'b10010010100100: data = 6'b010101;
12'b10010010100101: data = 6'b010101;
12'b10010010100110: data = 6'b010101;
12'b10010010100111: data = 6'b010101;
12'b10010010101000: data = 6'b010101;
12'b10010010101001: data = 6'b010101;
12'b10010010101010: data = 6'b010101;
12'b100101000000: data = 6'b010101;
12'b100101000001: data = 6'b010101;
12'b100101000010: data = 6'b010101;
12'b100101000011: data = 6'b010101;
12'b100101000100: data = 6'b010101;
12'b100101000101: data = 6'b010101;
12'b100101000110: data = 6'b010101;
12'b100101000111: data = 6'b010101;
12'b100101001000: data = 6'b010101;
12'b100101001001: data = 6'b010101;
12'b100101001010: data = 6'b010101;
12'b100101001011: data = 6'b010101;
12'b100101001100: data = 6'b010101;
12'b100101001101: data = 6'b010101;
12'b100101001110: data = 6'b010101;
12'b100101001111: data = 6'b010101;
12'b100101010000: data = 6'b010101;
12'b100101010001: data = 6'b010101;
12'b100101010010: data = 6'b010101;
12'b100101010011: data = 6'b010101;
12'b100101010100: data = 6'b010101;
12'b100101010101: data = 6'b010101;
12'b100101010110: data = 6'b010101;
12'b100101010111: data = 6'b010101;
12'b100101011000: data = 6'b010101;
12'b100101011001: data = 6'b101010;
12'b100101011010: data = 6'b101010;
12'b100101011011: data = 6'b101010;
12'b100101011100: data = 6'b010101;
12'b100101011101: data = 6'b000000;
12'b100101011110: data = 6'b000000;
12'b100101011111: data = 6'b010101;
12'b100101100000: data = 6'b010101;
12'b100101100001: data = 6'b010101;
12'b100101100010: data = 6'b010101;
12'b100101100011: data = 6'b101001;
12'b100101100100: data = 6'b101010;
12'b100101100101: data = 6'b101010;
12'b100101100110: data = 6'b101010;
12'b100101100111: data = 6'b101010;
12'b100101101000: data = 6'b101010;
12'b100101101001: data = 6'b101010;
12'b100101101010: data = 6'b101010;
12'b100101101011: data = 6'b101010;
12'b100101101100: data = 6'b101010;
12'b100101101101: data = 6'b101010;
12'b100101101110: data = 6'b101010;
12'b100101101111: data = 6'b101010;
12'b100101110000: data = 6'b101010;
12'b100101110001: data = 6'b101010;
12'b100101110010: data = 6'b101010;
12'b100101110011: data = 6'b101010;
12'b100101110100: data = 6'b101010;
12'b100101110101: data = 6'b101010;
12'b100101110110: data = 6'b101010;
12'b100101110111: data = 6'b101010;
12'b100101111000: data = 6'b101010;
12'b100101111001: data = 6'b101010;
12'b100101111010: data = 6'b101010;
12'b100101111011: data = 6'b101010;
12'b100101111100: data = 6'b111010;
12'b100101111101: data = 6'b111010;
12'b100101111110: data = 6'b111010;
12'b100101111111: data = 6'b111010;
12'b1001011000000: data = 6'b111010;
12'b1001011000001: data = 6'b101010;
12'b1001011000010: data = 6'b101010;
12'b1001011000011: data = 6'b101010;
12'b1001011000100: data = 6'b101010;
12'b1001011000101: data = 6'b101010;
12'b1001011000110: data = 6'b101010;
12'b1001011000111: data = 6'b101010;
12'b1001011001000: data = 6'b101010;
12'b1001011001001: data = 6'b101010;
12'b1001011001010: data = 6'b101010;
12'b1001011001011: data = 6'b101010;
12'b1001011001100: data = 6'b101010;
12'b1001011001101: data = 6'b101010;
12'b1001011001110: data = 6'b101010;
12'b1001011001111: data = 6'b101010;
12'b1001011010000: data = 6'b101010;
12'b1001011010001: data = 6'b101010;
12'b1001011010010: data = 6'b101010;
12'b1001011010011: data = 6'b101010;
12'b1001011010100: data = 6'b101010;
12'b1001011010101: data = 6'b101010;
12'b1001011010110: data = 6'b101010;
12'b1001011010111: data = 6'b101010;
12'b1001011011000: data = 6'b101010;
12'b1001011011001: data = 6'b101010;
12'b1001011011010: data = 6'b101010;
12'b1001011011011: data = 6'b101010;
12'b1001011011100: data = 6'b101010;
12'b1001011011101: data = 6'b101010;
12'b1001011011110: data = 6'b101010;
12'b1001011011111: data = 6'b101010;
12'b1001011100000: data = 6'b101010;
12'b1001011100001: data = 6'b101010;
12'b1001011100010: data = 6'b101010;
12'b1001011100011: data = 6'b101010;
12'b1001011100100: data = 6'b101010;
12'b1001011100101: data = 6'b101010;
12'b1001011100110: data = 6'b101010;
12'b1001011100111: data = 6'b101010;
12'b1001011101000: data = 6'b101010;
12'b1001011101001: data = 6'b101010;
12'b1001011101010: data = 6'b101010;
12'b1001011101011: data = 6'b101010;
12'b1001011101100: data = 6'b101010;
12'b1001011101101: data = 6'b101010;
12'b1001011101110: data = 6'b101010;
12'b1001011101111: data = 6'b101010;
12'b1001011110000: data = 6'b101010;
12'b1001011110001: data = 6'b101010;
12'b1001011110010: data = 6'b101010;
12'b1001011110011: data = 6'b101010;
12'b1001011110100: data = 6'b101010;
12'b1001011110101: data = 6'b101010;
12'b1001011110110: data = 6'b101010;
12'b1001011110111: data = 6'b101010;
12'b1001011111000: data = 6'b101010;
12'b1001011111001: data = 6'b101010;
12'b1001011111010: data = 6'b101010;
12'b1001011111011: data = 6'b101010;
12'b1001011111100: data = 6'b101010;
12'b1001011111101: data = 6'b101010;
12'b1001011111110: data = 6'b101010;
12'b1001011111111: data = 6'b101010;
12'b10010110000000: data = 6'b101010;
12'b10010110000001: data = 6'b101010;
12'b10010110000010: data = 6'b101010;
12'b10010110000011: data = 6'b101010;
12'b10010110000100: data = 6'b101010;
12'b10010110000101: data = 6'b101010;
12'b10010110000110: data = 6'b101001;
12'b10010110000111: data = 6'b010101;
12'b10010110001000: data = 6'b010101;
12'b10010110001001: data = 6'b010101;
12'b10010110001010: data = 6'b010101;
12'b10010110001011: data = 6'b010101;
12'b10010110001100: data = 6'b000000;
12'b10010110001101: data = 6'b000000;
12'b10010110001110: data = 6'b101010;
12'b10010110001111: data = 6'b101010;
12'b10010110010000: data = 6'b101010;
12'b10010110010001: data = 6'b101010;
12'b10010110010010: data = 6'b010101;
12'b10010110010011: data = 6'b010101;
12'b10010110010100: data = 6'b010101;
12'b10010110010101: data = 6'b010101;
12'b10010110010110: data = 6'b010101;
12'b10010110010111: data = 6'b010101;
12'b10010110011000: data = 6'b010101;
12'b10010110011001: data = 6'b010101;
12'b10010110011010: data = 6'b010101;
12'b10010110011011: data = 6'b010101;
12'b10010110011100: data = 6'b010101;
12'b10010110011101: data = 6'b010101;
12'b10010110011110: data = 6'b010101;
12'b10010110011111: data = 6'b010101;
12'b10010110100000: data = 6'b010101;
12'b10010110100001: data = 6'b010101;
12'b10010110100010: data = 6'b010101;
12'b10010110100011: data = 6'b010101;
12'b10010110100100: data = 6'b010101;
12'b10010110100101: data = 6'b010101;
12'b10010110100110: data = 6'b010101;
12'b10010110100111: data = 6'b010101;
12'b10010110101000: data = 6'b010101;
12'b10010110101001: data = 6'b010101;
12'b10010110101010: data = 6'b010101;
12'b100110000000: data = 6'b010101;
12'b100110000001: data = 6'b010101;
12'b100110000010: data = 6'b010101;
12'b100110000011: data = 6'b010101;
12'b100110000100: data = 6'b010101;
12'b100110000101: data = 6'b010101;
12'b100110000110: data = 6'b010101;
12'b100110000111: data = 6'b010101;
12'b100110001000: data = 6'b010101;
12'b100110001001: data = 6'b010101;
12'b100110001010: data = 6'b010101;
12'b100110001011: data = 6'b010101;
12'b100110001100: data = 6'b010101;
12'b100110001101: data = 6'b010101;
12'b100110001110: data = 6'b010101;
12'b100110001111: data = 6'b010101;
12'b100110010000: data = 6'b010101;
12'b100110010001: data = 6'b010101;
12'b100110010010: data = 6'b010101;
12'b100110010011: data = 6'b010101;
12'b100110010100: data = 6'b010101;
12'b100110010101: data = 6'b010101;
12'b100110010110: data = 6'b010101;
12'b100110010111: data = 6'b010101;
12'b100110011000: data = 6'b010101;
12'b100110011001: data = 6'b101010;
12'b100110011010: data = 6'b101010;
12'b100110011011: data = 6'b101010;
12'b100110011100: data = 6'b010101;
12'b100110011101: data = 6'b000000;
12'b100110011110: data = 6'b000000;
12'b100110011111: data = 6'b010101;
12'b100110100000: data = 6'b010101;
12'b100110100001: data = 6'b010101;
12'b100110100010: data = 6'b101001;
12'b100110100011: data = 6'b101010;
12'b100110100100: data = 6'b101010;
12'b100110100101: data = 6'b101010;
12'b100110100110: data = 6'b101010;
12'b100110100111: data = 6'b101010;
12'b100110101000: data = 6'b101010;
12'b100110101001: data = 6'b101010;
12'b100110101010: data = 6'b101010;
12'b100110101011: data = 6'b101010;
12'b100110101100: data = 6'b101010;
12'b100110101101: data = 6'b101010;
12'b100110101110: data = 6'b101010;
12'b100110101111: data = 6'b101010;
12'b100110110000: data = 6'b101010;
12'b100110110001: data = 6'b101010;
12'b100110110010: data = 6'b101010;
12'b100110110011: data = 6'b101010;
12'b100110110100: data = 6'b101010;
12'b100110110101: data = 6'b101010;
12'b100110110110: data = 6'b101010;
12'b100110110111: data = 6'b101010;
12'b100110111000: data = 6'b101010;
12'b100110111001: data = 6'b101010;
12'b100110111010: data = 6'b101010;
12'b100110111011: data = 6'b101010;
12'b100110111100: data = 6'b101010;
12'b100110111101: data = 6'b101010;
12'b100110111110: data = 6'b101010;
12'b100110111111: data = 6'b101010;
12'b1001101000000: data = 6'b101010;
12'b1001101000001: data = 6'b101010;
12'b1001101000010: data = 6'b101010;
12'b1001101000011: data = 6'b101010;
12'b1001101000100: data = 6'b101010;
12'b1001101000101: data = 6'b101010;
12'b1001101000110: data = 6'b101010;
12'b1001101000111: data = 6'b101010;
12'b1001101001000: data = 6'b101010;
12'b1001101001001: data = 6'b101010;
12'b1001101001010: data = 6'b101010;
12'b1001101001011: data = 6'b101010;
12'b1001101001100: data = 6'b101010;
12'b1001101001101: data = 6'b101010;
12'b1001101001110: data = 6'b101010;
12'b1001101001111: data = 6'b101010;
12'b1001101010000: data = 6'b101010;
12'b1001101010001: data = 6'b101010;
12'b1001101010010: data = 6'b101010;
12'b1001101010011: data = 6'b101010;
12'b1001101010100: data = 6'b101010;
12'b1001101010101: data = 6'b101010;
12'b1001101010110: data = 6'b101010;
12'b1001101010111: data = 6'b101010;
12'b1001101011000: data = 6'b101010;
12'b1001101011001: data = 6'b101010;
12'b1001101011010: data = 6'b101010;
12'b1001101011011: data = 6'b101010;
12'b1001101011100: data = 6'b101010;
12'b1001101011101: data = 6'b101010;
12'b1001101011110: data = 6'b101010;
12'b1001101011111: data = 6'b101010;
12'b1001101100000: data = 6'b101010;
12'b1001101100001: data = 6'b101010;
12'b1001101100010: data = 6'b101010;
12'b1001101100011: data = 6'b101010;
12'b1001101100100: data = 6'b101010;
12'b1001101100101: data = 6'b101010;
12'b1001101100110: data = 6'b101010;
12'b1001101100111: data = 6'b101010;
12'b1001101101000: data = 6'b101010;
12'b1001101101001: data = 6'b101010;
12'b1001101101010: data = 6'b101010;
12'b1001101101011: data = 6'b101010;
12'b1001101101100: data = 6'b101010;
12'b1001101101101: data = 6'b101010;
12'b1001101101110: data = 6'b101010;
12'b1001101101111: data = 6'b101010;
12'b1001101110000: data = 6'b101010;
12'b1001101110001: data = 6'b101010;
12'b1001101110010: data = 6'b101010;
12'b1001101110011: data = 6'b101010;
12'b1001101110100: data = 6'b101010;
12'b1001101110101: data = 6'b101010;
12'b1001101110110: data = 6'b101010;
12'b1001101110111: data = 6'b101010;
12'b1001101111000: data = 6'b101010;
12'b1001101111001: data = 6'b101010;
12'b1001101111010: data = 6'b101010;
12'b1001101111011: data = 6'b101010;
12'b1001101111100: data = 6'b101010;
12'b1001101111101: data = 6'b101010;
12'b1001101111110: data = 6'b101010;
12'b1001101111111: data = 6'b101010;
12'b10011010000000: data = 6'b101010;
12'b10011010000001: data = 6'b101010;
12'b10011010000010: data = 6'b101010;
12'b10011010000011: data = 6'b101010;
12'b10011010000100: data = 6'b101010;
12'b10011010000101: data = 6'b101010;
12'b10011010000110: data = 6'b101010;
12'b10011010000111: data = 6'b101010;
12'b10011010001000: data = 6'b101001;
12'b10011010001001: data = 6'b010101;
12'b10011010001010: data = 6'b010101;
12'b10011010001011: data = 6'b010101;
12'b10011010001100: data = 6'b000000;
12'b10011010001101: data = 6'b000000;
12'b10011010001110: data = 6'b101010;
12'b10011010001111: data = 6'b101010;
12'b10011010010000: data = 6'b101010;
12'b10011010010001: data = 6'b101010;
12'b10011010010010: data = 6'b010101;
12'b10011010010011: data = 6'b010101;
12'b10011010010100: data = 6'b010101;
12'b10011010010101: data = 6'b010101;
12'b10011010010110: data = 6'b010101;
12'b10011010010111: data = 6'b010101;
12'b10011010011000: data = 6'b010101;
12'b10011010011001: data = 6'b010101;
12'b10011010011010: data = 6'b010101;
12'b10011010011011: data = 6'b010101;
12'b10011010011100: data = 6'b010101;
12'b10011010011101: data = 6'b010101;
12'b10011010011110: data = 6'b010101;
12'b10011010011111: data = 6'b010101;
12'b10011010100000: data = 6'b010101;
12'b10011010100001: data = 6'b010101;
12'b10011010100010: data = 6'b010101;
12'b10011010100011: data = 6'b010101;
12'b10011010100100: data = 6'b010101;
12'b10011010100101: data = 6'b010101;
12'b10011010100110: data = 6'b010101;
12'b10011010100111: data = 6'b010101;
12'b10011010101000: data = 6'b010101;
12'b10011010101001: data = 6'b010101;
12'b10011010101010: data = 6'b010101;
12'b100111000000: data = 6'b010101;
12'b100111000001: data = 6'b010101;
12'b100111000010: data = 6'b010101;
12'b100111000011: data = 6'b010101;
12'b100111000100: data = 6'b010101;
12'b100111000101: data = 6'b010101;
12'b100111000110: data = 6'b010101;
12'b100111000111: data = 6'b010101;
12'b100111001000: data = 6'b010101;
12'b100111001001: data = 6'b010101;
12'b100111001010: data = 6'b010101;
12'b100111001011: data = 6'b010101;
12'b100111001100: data = 6'b010101;
12'b100111001101: data = 6'b010101;
12'b100111001110: data = 6'b010101;
12'b100111001111: data = 6'b010101;
12'b100111010000: data = 6'b010101;
12'b100111010001: data = 6'b010101;
12'b100111010010: data = 6'b010101;
12'b100111010011: data = 6'b010101;
12'b100111010100: data = 6'b010101;
12'b100111010101: data = 6'b010101;
12'b100111010110: data = 6'b010101;
12'b100111010111: data = 6'b010101;
12'b100111011000: data = 6'b010101;
12'b100111011001: data = 6'b101010;
12'b100111011010: data = 6'b101010;
12'b100111011011: data = 6'b101010;
12'b100111011100: data = 6'b010101;
12'b100111011101: data = 6'b000000;
12'b100111011110: data = 6'b000000;
12'b100111011111: data = 6'b010101;
12'b100111100000: data = 6'b010101;
12'b100111100001: data = 6'b010101;
12'b100111100010: data = 6'b101001;
12'b100111100011: data = 6'b101010;
12'b100111100100: data = 6'b101010;
12'b100111100101: data = 6'b101010;
12'b100111100110: data = 6'b101010;
12'b100111100111: data = 6'b101010;
12'b100111101000: data = 6'b101010;
12'b100111101001: data = 6'b101010;
12'b100111101010: data = 6'b101010;
12'b100111101011: data = 6'b101010;
12'b100111101100: data = 6'b101010;
12'b100111101101: data = 6'b101010;
12'b100111101110: data = 6'b101010;
12'b100111101111: data = 6'b101010;
12'b100111110000: data = 6'b101010;
12'b100111110001: data = 6'b101010;
12'b100111110010: data = 6'b101010;
12'b100111110011: data = 6'b101010;
12'b100111110100: data = 6'b101010;
12'b100111110101: data = 6'b101010;
12'b100111110110: data = 6'b101010;
12'b100111110111: data = 6'b101010;
12'b100111111000: data = 6'b101010;
12'b100111111001: data = 6'b101010;
12'b100111111010: data = 6'b101010;
12'b100111111011: data = 6'b101010;
12'b100111111100: data = 6'b101010;
12'b100111111101: data = 6'b101010;
12'b100111111110: data = 6'b101010;
12'b100111111111: data = 6'b101010;
12'b1001111000000: data = 6'b101010;
12'b1001111000001: data = 6'b101010;
12'b1001111000010: data = 6'b101010;
12'b1001111000011: data = 6'b101010;
12'b1001111000100: data = 6'b101010;
12'b1001111000101: data = 6'b101010;
12'b1001111000110: data = 6'b101010;
12'b1001111000111: data = 6'b101010;
12'b1001111001000: data = 6'b101010;
12'b1001111001001: data = 6'b101010;
12'b1001111001010: data = 6'b101010;
12'b1001111001011: data = 6'b101010;
12'b1001111001100: data = 6'b101010;
12'b1001111001101: data = 6'b101010;
12'b1001111001110: data = 6'b101010;
12'b1001111001111: data = 6'b101010;
12'b1001111010000: data = 6'b101010;
12'b1001111010001: data = 6'b101010;
12'b1001111010010: data = 6'b101010;
12'b1001111010011: data = 6'b101010;
12'b1001111010100: data = 6'b101010;
12'b1001111010101: data = 6'b101010;
12'b1001111010110: data = 6'b101010;
12'b1001111010111: data = 6'b101010;
12'b1001111011000: data = 6'b101010;
12'b1001111011001: data = 6'b101010;
12'b1001111011010: data = 6'b101010;
12'b1001111011011: data = 6'b101010;
12'b1001111011100: data = 6'b101010;
12'b1001111011101: data = 6'b101010;
12'b1001111011110: data = 6'b101010;
12'b1001111011111: data = 6'b101010;
12'b1001111100000: data = 6'b101010;
12'b1001111100001: data = 6'b101010;
12'b1001111100010: data = 6'b101010;
12'b1001111100011: data = 6'b101010;
12'b1001111100100: data = 6'b101010;
12'b1001111100101: data = 6'b101010;
12'b1001111100110: data = 6'b101010;
12'b1001111100111: data = 6'b101010;
12'b1001111101000: data = 6'b101010;
12'b1001111101001: data = 6'b101010;
12'b1001111101010: data = 6'b101010;
12'b1001111101011: data = 6'b101010;
12'b1001111101100: data = 6'b101010;
12'b1001111101101: data = 6'b101010;
12'b1001111101110: data = 6'b101010;
12'b1001111101111: data = 6'b101010;
12'b1001111110000: data = 6'b101010;
12'b1001111110001: data = 6'b101010;
12'b1001111110010: data = 6'b101010;
12'b1001111110011: data = 6'b101010;
12'b1001111110100: data = 6'b101010;
12'b1001111110101: data = 6'b101010;
12'b1001111110110: data = 6'b101010;
12'b1001111110111: data = 6'b101010;
12'b1001111111000: data = 6'b101010;
12'b1001111111001: data = 6'b101010;
12'b1001111111010: data = 6'b101010;
12'b1001111111011: data = 6'b101010;
12'b1001111111100: data = 6'b101010;
12'b1001111111101: data = 6'b101010;
12'b1001111111110: data = 6'b101010;
12'b1001111111111: data = 6'b101010;
12'b10011110000000: data = 6'b101010;
12'b10011110000001: data = 6'b101010;
12'b10011110000010: data = 6'b101010;
12'b10011110000011: data = 6'b101010;
12'b10011110000100: data = 6'b101010;
12'b10011110000101: data = 6'b101010;
12'b10011110000110: data = 6'b101010;
12'b10011110000111: data = 6'b101010;
12'b10011110001000: data = 6'b101001;
12'b10011110001001: data = 6'b010101;
12'b10011110001010: data = 6'b010101;
12'b10011110001011: data = 6'b010101;
12'b10011110001100: data = 6'b000000;
12'b10011110001101: data = 6'b000000;
12'b10011110001110: data = 6'b101010;
12'b10011110001111: data = 6'b101010;
12'b10011110010000: data = 6'b101010;
12'b10011110010001: data = 6'b101010;
12'b10011110010010: data = 6'b010101;
12'b10011110010011: data = 6'b010101;
12'b10011110010100: data = 6'b010101;
12'b10011110010101: data = 6'b010101;
12'b10011110010110: data = 6'b010101;
12'b10011110010111: data = 6'b010101;
12'b10011110011000: data = 6'b010101;
12'b10011110011001: data = 6'b010101;
12'b10011110011010: data = 6'b010101;
12'b10011110011011: data = 6'b010101;
12'b10011110011100: data = 6'b010101;
12'b10011110011101: data = 6'b010101;
12'b10011110011110: data = 6'b010101;
12'b10011110011111: data = 6'b010101;
12'b10011110100000: data = 6'b010101;
12'b10011110100001: data = 6'b010101;
12'b10011110100010: data = 6'b010101;
12'b10011110100011: data = 6'b010101;
12'b10011110100100: data = 6'b010101;
12'b10011110100101: data = 6'b010101;
12'b10011110100110: data = 6'b010101;
12'b10011110100111: data = 6'b010101;
12'b10011110101000: data = 6'b010101;
12'b10011110101001: data = 6'b010101;
12'b10011110101010: data = 6'b010101;
12'b101000000000: data = 6'b010101;
12'b101000000001: data = 6'b010101;
12'b101000000010: data = 6'b010101;
12'b101000000011: data = 6'b010101;
12'b101000000100: data = 6'b010101;
12'b101000000101: data = 6'b010101;
12'b101000000110: data = 6'b010101;
12'b101000000111: data = 6'b010101;
12'b101000001000: data = 6'b010101;
12'b101000001001: data = 6'b010101;
12'b101000001010: data = 6'b010101;
12'b101000001011: data = 6'b010101;
12'b101000001100: data = 6'b010101;
12'b101000001101: data = 6'b010101;
12'b101000001110: data = 6'b010101;
12'b101000001111: data = 6'b010101;
12'b101000010000: data = 6'b010101;
12'b101000010001: data = 6'b010101;
12'b101000010010: data = 6'b010101;
12'b101000010011: data = 6'b010101;
12'b101000010100: data = 6'b010101;
12'b101000010101: data = 6'b010101;
12'b101000010110: data = 6'b010101;
12'b101000010111: data = 6'b010101;
12'b101000011000: data = 6'b010101;
12'b101000011001: data = 6'b101010;
12'b101000011010: data = 6'b101010;
12'b101000011011: data = 6'b101010;
12'b101000011100: data = 6'b010101;
12'b101000011101: data = 6'b000000;
12'b101000011110: data = 6'b000000;
12'b101000011111: data = 6'b010101;
12'b101000100000: data = 6'b010101;
12'b101000100001: data = 6'b010101;
12'b101000100010: data = 6'b101010;
12'b101000100011: data = 6'b101010;
12'b101000100100: data = 6'b101010;
12'b101000100101: data = 6'b101010;
12'b101000100110: data = 6'b101010;
12'b101000100111: data = 6'b101010;
12'b101000101000: data = 6'b101010;
12'b101000101001: data = 6'b101010;
12'b101000101010: data = 6'b101010;
12'b101000101011: data = 6'b101010;
12'b101000101100: data = 6'b101010;
12'b101000101101: data = 6'b101010;
12'b101000101110: data = 6'b101010;
12'b101000101111: data = 6'b101010;
12'b101000110000: data = 6'b101010;
12'b101000110001: data = 6'b101010;
12'b101000110010: data = 6'b101010;
12'b101000110011: data = 6'b101010;
12'b101000110100: data = 6'b101010;
12'b101000110101: data = 6'b101010;
12'b101000110110: data = 6'b101010;
12'b101000110111: data = 6'b101010;
12'b101000111000: data = 6'b101010;
12'b101000111001: data = 6'b101010;
12'b101000111010: data = 6'b101010;
12'b101000111011: data = 6'b101010;
12'b101000111100: data = 6'b101010;
12'b101000111101: data = 6'b101010;
12'b101000111110: data = 6'b101010;
12'b101000111111: data = 6'b101010;
12'b1010001000000: data = 6'b101010;
12'b1010001000001: data = 6'b101010;
12'b1010001000010: data = 6'b101010;
12'b1010001000011: data = 6'b101010;
12'b1010001000100: data = 6'b101010;
12'b1010001000101: data = 6'b101010;
12'b1010001000110: data = 6'b101010;
12'b1010001000111: data = 6'b101010;
12'b1010001001000: data = 6'b101010;
12'b1010001001001: data = 6'b101010;
12'b1010001001010: data = 6'b101010;
12'b1010001001011: data = 6'b101010;
12'b1010001001100: data = 6'b101010;
12'b1010001001101: data = 6'b101010;
12'b1010001001110: data = 6'b101010;
12'b1010001001111: data = 6'b101010;
12'b1010001010000: data = 6'b101010;
12'b1010001010001: data = 6'b101010;
12'b1010001010010: data = 6'b101010;
12'b1010001010011: data = 6'b101010;
12'b1010001010100: data = 6'b101010;
12'b1010001010101: data = 6'b101010;
12'b1010001010110: data = 6'b101010;
12'b1010001010111: data = 6'b101010;
12'b1010001011000: data = 6'b101010;
12'b1010001011001: data = 6'b101010;
12'b1010001011010: data = 6'b101010;
12'b1010001011011: data = 6'b101010;
12'b1010001011100: data = 6'b101010;
12'b1010001011101: data = 6'b101010;
12'b1010001011110: data = 6'b101010;
12'b1010001011111: data = 6'b101010;
12'b1010001100000: data = 6'b101010;
12'b1010001100001: data = 6'b101010;
12'b1010001100010: data = 6'b101010;
12'b1010001100011: data = 6'b101010;
12'b1010001100100: data = 6'b101010;
12'b1010001100101: data = 6'b101010;
12'b1010001100110: data = 6'b101010;
12'b1010001100111: data = 6'b101010;
12'b1010001101000: data = 6'b101010;
12'b1010001101001: data = 6'b101010;
12'b1010001101010: data = 6'b101010;
12'b1010001101011: data = 6'b101010;
12'b1010001101100: data = 6'b101010;
12'b1010001101101: data = 6'b101010;
12'b1010001101110: data = 6'b101010;
12'b1010001101111: data = 6'b101010;
12'b1010001110000: data = 6'b101010;
12'b1010001110001: data = 6'b101010;
12'b1010001110010: data = 6'b101010;
12'b1010001110011: data = 6'b101010;
12'b1010001110100: data = 6'b101010;
12'b1010001110101: data = 6'b101010;
12'b1010001110110: data = 6'b101010;
12'b1010001110111: data = 6'b101010;
12'b1010001111000: data = 6'b101010;
12'b1010001111001: data = 6'b101010;
12'b1010001111010: data = 6'b101010;
12'b1010001111011: data = 6'b101010;
12'b1010001111100: data = 6'b101010;
12'b1010001111101: data = 6'b101010;
12'b1010001111110: data = 6'b101010;
12'b1010001111111: data = 6'b101010;
12'b10100010000000: data = 6'b101010;
12'b10100010000001: data = 6'b101010;
12'b10100010000010: data = 6'b101010;
12'b10100010000011: data = 6'b101010;
12'b10100010000100: data = 6'b101010;
12'b10100010000101: data = 6'b101010;
12'b10100010000110: data = 6'b101010;
12'b10100010000111: data = 6'b101010;
12'b10100010001000: data = 6'b101001;
12'b10100010001001: data = 6'b010101;
12'b10100010001010: data = 6'b010101;
12'b10100010001011: data = 6'b010101;
12'b10100010001100: data = 6'b000000;
12'b10100010001101: data = 6'b000000;
12'b10100010001110: data = 6'b101010;
12'b10100010001111: data = 6'b101010;
12'b10100010010000: data = 6'b101010;
12'b10100010010001: data = 6'b101010;
12'b10100010010010: data = 6'b010101;
12'b10100010010011: data = 6'b010101;
12'b10100010010100: data = 6'b010101;
12'b10100010010101: data = 6'b010101;
12'b10100010010110: data = 6'b010101;
12'b10100010010111: data = 6'b010101;
12'b10100010011000: data = 6'b010101;
12'b10100010011001: data = 6'b010101;
12'b10100010011010: data = 6'b010101;
12'b10100010011011: data = 6'b010101;
12'b10100010011100: data = 6'b010101;
12'b10100010011101: data = 6'b010101;
12'b10100010011110: data = 6'b010101;
12'b10100010011111: data = 6'b010101;
12'b10100010100000: data = 6'b010101;
12'b10100010100001: data = 6'b010101;
12'b10100010100010: data = 6'b010101;
12'b10100010100011: data = 6'b010101;
12'b10100010100100: data = 6'b010101;
12'b10100010100101: data = 6'b010101;
12'b10100010100110: data = 6'b010101;
12'b10100010100111: data = 6'b010101;
12'b10100010101000: data = 6'b010101;
12'b10100010101001: data = 6'b010101;
12'b10100010101010: data = 6'b010101;
12'b101001000000: data = 6'b010101;
12'b101001000001: data = 6'b010101;
12'b101001000010: data = 6'b010101;
12'b101001000011: data = 6'b010101;
12'b101001000100: data = 6'b010101;
12'b101001000101: data = 6'b010101;
12'b101001000110: data = 6'b010101;
12'b101001000111: data = 6'b010101;
12'b101001001000: data = 6'b010101;
12'b101001001001: data = 6'b010101;
12'b101001001010: data = 6'b010101;
12'b101001001011: data = 6'b010101;
12'b101001001100: data = 6'b010101;
12'b101001001101: data = 6'b010101;
12'b101001001110: data = 6'b010101;
12'b101001001111: data = 6'b010101;
12'b101001010000: data = 6'b010101;
12'b101001010001: data = 6'b010101;
12'b101001010010: data = 6'b010101;
12'b101001010011: data = 6'b010101;
12'b101001010100: data = 6'b010101;
12'b101001010101: data = 6'b010101;
12'b101001010110: data = 6'b010101;
12'b101001010111: data = 6'b010101;
12'b101001011000: data = 6'b010101;
12'b101001011001: data = 6'b101010;
12'b101001011010: data = 6'b101010;
12'b101001011011: data = 6'b101010;
12'b101001011100: data = 6'b010101;
12'b101001011101: data = 6'b000000;
12'b101001011110: data = 6'b000000;
12'b101001011111: data = 6'b010101;
12'b101001100000: data = 6'b010101;
12'b101001100001: data = 6'b010101;
12'b101001100010: data = 6'b101010;
12'b101001100011: data = 6'b101010;
12'b101001100100: data = 6'b101010;
12'b101001100101: data = 6'b101010;
12'b101001100110: data = 6'b101010;
12'b101001100111: data = 6'b101010;
12'b101001101000: data = 6'b101010;
12'b101001101001: data = 6'b101010;
12'b101001101010: data = 6'b101010;
12'b101001101011: data = 6'b101010;
12'b101001101100: data = 6'b101010;
12'b101001101101: data = 6'b101010;
12'b101001101110: data = 6'b101010;
12'b101001101111: data = 6'b101010;
12'b101001110000: data = 6'b101010;
12'b101001110001: data = 6'b101010;
12'b101001110010: data = 6'b101010;
12'b101001110011: data = 6'b101010;
12'b101001110100: data = 6'b101010;
12'b101001110101: data = 6'b101010;
12'b101001110110: data = 6'b101010;
12'b101001110111: data = 6'b101010;
12'b101001111000: data = 6'b101010;
12'b101001111001: data = 6'b101010;
12'b101001111010: data = 6'b101010;
12'b101001111011: data = 6'b101010;
12'b101001111100: data = 6'b101010;
12'b101001111101: data = 6'b101010;
12'b101001111110: data = 6'b101010;
12'b101001111111: data = 6'b101010;
12'b1010011000000: data = 6'b101010;
12'b1010011000001: data = 6'b101010;
12'b1010011000010: data = 6'b101010;
12'b1010011000011: data = 6'b101010;
12'b1010011000100: data = 6'b101010;
12'b1010011000101: data = 6'b101010;
12'b1010011000110: data = 6'b101010;
12'b1010011000111: data = 6'b101010;
12'b1010011001000: data = 6'b101010;
12'b1010011001001: data = 6'b101010;
12'b1010011001010: data = 6'b101010;
12'b1010011001011: data = 6'b101010;
12'b1010011001100: data = 6'b101010;
12'b1010011001101: data = 6'b101010;
12'b1010011001110: data = 6'b101010;
12'b1010011001111: data = 6'b101010;
12'b1010011010000: data = 6'b101010;
12'b1010011010001: data = 6'b101010;
12'b1010011010010: data = 6'b101010;
12'b1010011010011: data = 6'b101010;
12'b1010011010100: data = 6'b101010;
12'b1010011010101: data = 6'b101010;
12'b1010011010110: data = 6'b101010;
12'b1010011010111: data = 6'b101010;
12'b1010011011000: data = 6'b101010;
12'b1010011011001: data = 6'b101010;
12'b1010011011010: data = 6'b101010;
12'b1010011011011: data = 6'b101010;
12'b1010011011100: data = 6'b101010;
12'b1010011011101: data = 6'b101010;
12'b1010011011110: data = 6'b101010;
12'b1010011011111: data = 6'b101010;
12'b1010011100000: data = 6'b101010;
12'b1010011100001: data = 6'b101010;
12'b1010011100010: data = 6'b101010;
12'b1010011100011: data = 6'b101010;
12'b1010011100100: data = 6'b101010;
12'b1010011100101: data = 6'b101010;
12'b1010011100110: data = 6'b101010;
12'b1010011100111: data = 6'b101010;
12'b1010011101000: data = 6'b101010;
12'b1010011101001: data = 6'b101010;
12'b1010011101010: data = 6'b101010;
12'b1010011101011: data = 6'b101010;
12'b1010011101100: data = 6'b101010;
12'b1010011101101: data = 6'b101010;
12'b1010011101110: data = 6'b101010;
12'b1010011101111: data = 6'b101010;
12'b1010011110000: data = 6'b101010;
12'b1010011110001: data = 6'b101010;
12'b1010011110010: data = 6'b101010;
12'b1010011110011: data = 6'b101010;
12'b1010011110100: data = 6'b101010;
12'b1010011110101: data = 6'b101010;
12'b1010011110110: data = 6'b101010;
12'b1010011110111: data = 6'b101010;
12'b1010011111000: data = 6'b101010;
12'b1010011111001: data = 6'b101010;
12'b1010011111010: data = 6'b101010;
12'b1010011111011: data = 6'b101010;
12'b1010011111100: data = 6'b101010;
12'b1010011111101: data = 6'b101010;
12'b1010011111110: data = 6'b101010;
12'b1010011111111: data = 6'b101010;
12'b10100110000000: data = 6'b101010;
12'b10100110000001: data = 6'b101010;
12'b10100110000010: data = 6'b101010;
12'b10100110000011: data = 6'b101010;
12'b10100110000100: data = 6'b101010;
12'b10100110000101: data = 6'b101010;
12'b10100110000110: data = 6'b101010;
12'b10100110000111: data = 6'b101010;
12'b10100110001000: data = 6'b101010;
12'b10100110001001: data = 6'b010101;
12'b10100110001010: data = 6'b010101;
12'b10100110001011: data = 6'b010101;
12'b10100110001100: data = 6'b000000;
12'b10100110001101: data = 6'b000000;
12'b10100110001110: data = 6'b101010;
12'b10100110001111: data = 6'b101010;
12'b10100110010000: data = 6'b101010;
12'b10100110010001: data = 6'b101010;
12'b10100110010010: data = 6'b010101;
12'b10100110010011: data = 6'b010101;
12'b10100110010100: data = 6'b010101;
12'b10100110010101: data = 6'b010101;
12'b10100110010110: data = 6'b010101;
12'b10100110010111: data = 6'b010101;
12'b10100110011000: data = 6'b010101;
12'b10100110011001: data = 6'b010101;
12'b10100110011010: data = 6'b010101;
12'b10100110011011: data = 6'b010101;
12'b10100110011100: data = 6'b010101;
12'b10100110011101: data = 6'b010101;
12'b10100110011110: data = 6'b010101;
12'b10100110011111: data = 6'b010101;
12'b10100110100000: data = 6'b010101;
12'b10100110100001: data = 6'b010101;
12'b10100110100010: data = 6'b010101;
12'b10100110100011: data = 6'b010101;
12'b10100110100100: data = 6'b010101;
12'b10100110100101: data = 6'b010101;
12'b10100110100110: data = 6'b010101;
12'b10100110100111: data = 6'b010101;
12'b10100110101000: data = 6'b010101;
12'b10100110101001: data = 6'b010101;
12'b10100110101010: data = 6'b010101;
12'b101010000000: data = 6'b010101;
12'b101010000001: data = 6'b010101;
12'b101010000010: data = 6'b010101;
12'b101010000011: data = 6'b010101;
12'b101010000100: data = 6'b010101;
12'b101010000101: data = 6'b010101;
12'b101010000110: data = 6'b010101;
12'b101010000111: data = 6'b010101;
12'b101010001000: data = 6'b010101;
12'b101010001001: data = 6'b010101;
12'b101010001010: data = 6'b010101;
12'b101010001011: data = 6'b010101;
12'b101010001100: data = 6'b010101;
12'b101010001101: data = 6'b010101;
12'b101010001110: data = 6'b010101;
12'b101010001111: data = 6'b010101;
12'b101010010000: data = 6'b010101;
12'b101010010001: data = 6'b010101;
12'b101010010010: data = 6'b010101;
12'b101010010011: data = 6'b010101;
12'b101010010100: data = 6'b010101;
12'b101010010101: data = 6'b010101;
12'b101010010110: data = 6'b010101;
12'b101010010111: data = 6'b010101;
12'b101010011000: data = 6'b010101;
12'b101010011001: data = 6'b101010;
12'b101010011010: data = 6'b101010;
12'b101010011011: data = 6'b101010;
12'b101010011100: data = 6'b010101;
12'b101010011101: data = 6'b000000;
12'b101010011110: data = 6'b000000;
12'b101010011111: data = 6'b010101;
12'b101010100000: data = 6'b010101;
12'b101010100001: data = 6'b010101;
12'b101010100010: data = 6'b101010;
12'b101010100011: data = 6'b101010;
12'b101010100100: data = 6'b101010;
12'b101010100101: data = 6'b101010;
12'b101010100110: data = 6'b101010;
12'b101010100111: data = 6'b101010;
12'b101010101000: data = 6'b101010;
12'b101010101001: data = 6'b101010;
12'b101010101010: data = 6'b101010;
12'b101010101011: data = 6'b101010;
12'b101010101100: data = 6'b101010;
12'b101010101101: data = 6'b101010;
12'b101010101110: data = 6'b101010;
12'b101010101111: data = 6'b101010;
12'b101010110000: data = 6'b101010;
12'b101010110001: data = 6'b101010;
12'b101010110010: data = 6'b101010;
12'b101010110011: data = 6'b101010;
12'b101010110100: data = 6'b101010;
12'b101010110101: data = 6'b101010;
12'b101010110110: data = 6'b101010;
12'b101010110111: data = 6'b101010;
12'b101010111000: data = 6'b101010;
12'b101010111001: data = 6'b101010;
12'b101010111010: data = 6'b101010;
12'b101010111011: data = 6'b101010;
12'b101010111100: data = 6'b101010;
12'b101010111101: data = 6'b101010;
12'b101010111110: data = 6'b101010;
12'b101010111111: data = 6'b101010;
12'b1010101000000: data = 6'b101010;
12'b1010101000001: data = 6'b101010;
12'b1010101000010: data = 6'b101010;
12'b1010101000011: data = 6'b101010;
12'b1010101000100: data = 6'b101010;
12'b1010101000101: data = 6'b101010;
12'b1010101000110: data = 6'b101010;
12'b1010101000111: data = 6'b101010;
12'b1010101001000: data = 6'b101010;
12'b1010101001001: data = 6'b101010;
12'b1010101001010: data = 6'b101010;
12'b1010101001011: data = 6'b101010;
12'b1010101001100: data = 6'b101010;
12'b1010101001101: data = 6'b101010;
12'b1010101001110: data = 6'b101010;
12'b1010101001111: data = 6'b101010;
12'b1010101010000: data = 6'b101010;
12'b1010101010001: data = 6'b101010;
12'b1010101010010: data = 6'b101010;
12'b1010101010011: data = 6'b101010;
12'b1010101010100: data = 6'b101010;
12'b1010101010101: data = 6'b101010;
12'b1010101010110: data = 6'b101010;
12'b1010101010111: data = 6'b101010;
12'b1010101011000: data = 6'b101010;
12'b1010101011001: data = 6'b101010;
12'b1010101011010: data = 6'b101010;
12'b1010101011011: data = 6'b101010;
12'b1010101011100: data = 6'b101010;
12'b1010101011101: data = 6'b101010;
12'b1010101011110: data = 6'b101010;
12'b1010101011111: data = 6'b101010;
12'b1010101100000: data = 6'b101010;
12'b1010101100001: data = 6'b101010;
12'b1010101100010: data = 6'b101010;
12'b1010101100011: data = 6'b101010;
12'b1010101100100: data = 6'b101010;
12'b1010101100101: data = 6'b101010;
12'b1010101100110: data = 6'b101010;
12'b1010101100111: data = 6'b101010;
12'b1010101101000: data = 6'b101010;
12'b1010101101001: data = 6'b101010;
12'b1010101101010: data = 6'b101010;
12'b1010101101011: data = 6'b101010;
12'b1010101101100: data = 6'b101010;
12'b1010101101101: data = 6'b101010;
12'b1010101101110: data = 6'b101010;
12'b1010101101111: data = 6'b101010;
12'b1010101110000: data = 6'b101010;
12'b1010101110001: data = 6'b101010;
12'b1010101110010: data = 6'b101010;
12'b1010101110011: data = 6'b101010;
12'b1010101110100: data = 6'b101010;
12'b1010101110101: data = 6'b101010;
12'b1010101110110: data = 6'b101010;
12'b1010101110111: data = 6'b101010;
12'b1010101111000: data = 6'b101010;
12'b1010101111001: data = 6'b101010;
12'b1010101111010: data = 6'b101010;
12'b1010101111011: data = 6'b101010;
12'b1010101111100: data = 6'b101010;
12'b1010101111101: data = 6'b101010;
12'b1010101111110: data = 6'b101010;
12'b1010101111111: data = 6'b101010;
12'b10101010000000: data = 6'b101010;
12'b10101010000001: data = 6'b101010;
12'b10101010000010: data = 6'b101010;
12'b10101010000011: data = 6'b101010;
12'b10101010000100: data = 6'b101010;
12'b10101010000101: data = 6'b101010;
12'b10101010000110: data = 6'b101010;
12'b10101010000111: data = 6'b101010;
12'b10101010001000: data = 6'b101010;
12'b10101010001001: data = 6'b010101;
12'b10101010001010: data = 6'b010101;
12'b10101010001011: data = 6'b010101;
12'b10101010001100: data = 6'b000000;
12'b10101010001101: data = 6'b000000;
12'b10101010001110: data = 6'b101010;
12'b10101010001111: data = 6'b101010;
12'b10101010010000: data = 6'b101010;
12'b10101010010001: data = 6'b101010;
12'b10101010010010: data = 6'b010101;
12'b10101010010011: data = 6'b010101;
12'b10101010010100: data = 6'b010101;
12'b10101010010101: data = 6'b010101;
12'b10101010010110: data = 6'b010101;
12'b10101010010111: data = 6'b010101;
12'b10101010011000: data = 6'b010101;
12'b10101010011001: data = 6'b010101;
12'b10101010011010: data = 6'b010101;
12'b10101010011011: data = 6'b010101;
12'b10101010011100: data = 6'b010101;
12'b10101010011101: data = 6'b010101;
12'b10101010011110: data = 6'b010101;
12'b10101010011111: data = 6'b010101;
12'b10101010100000: data = 6'b010101;
12'b10101010100001: data = 6'b010101;
12'b10101010100010: data = 6'b010101;
12'b10101010100011: data = 6'b010101;
12'b10101010100100: data = 6'b010101;
12'b10101010100101: data = 6'b010101;
12'b10101010100110: data = 6'b010101;
12'b10101010100111: data = 6'b010101;
12'b10101010101000: data = 6'b010101;
12'b10101010101001: data = 6'b010101;
12'b10101010101010: data = 6'b010101;
12'b101011000000: data = 6'b010101;
12'b101011000001: data = 6'b010101;
12'b101011000010: data = 6'b010101;
12'b101011000011: data = 6'b010101;
12'b101011000100: data = 6'b010101;
12'b101011000101: data = 6'b010101;
12'b101011000110: data = 6'b010101;
12'b101011000111: data = 6'b010101;
12'b101011001000: data = 6'b010101;
12'b101011001001: data = 6'b010101;
12'b101011001010: data = 6'b010101;
12'b101011001011: data = 6'b010101;
12'b101011001100: data = 6'b010101;
12'b101011001101: data = 6'b010101;
12'b101011001110: data = 6'b010101;
12'b101011001111: data = 6'b010101;
12'b101011010000: data = 6'b010101;
12'b101011010001: data = 6'b010101;
12'b101011010010: data = 6'b010101;
12'b101011010011: data = 6'b010101;
12'b101011010100: data = 6'b010101;
12'b101011010101: data = 6'b010101;
12'b101011010110: data = 6'b010101;
12'b101011010111: data = 6'b010101;
12'b101011011000: data = 6'b010101;
12'b101011011001: data = 6'b101010;
12'b101011011010: data = 6'b101010;
12'b101011011011: data = 6'b101010;
12'b101011011100: data = 6'b010101;
12'b101011011101: data = 6'b000000;
12'b101011011110: data = 6'b000000;
12'b101011011111: data = 6'b010101;
12'b101011100000: data = 6'b010101;
12'b101011100001: data = 6'b010101;
12'b101011100010: data = 6'b101010;
12'b101011100011: data = 6'b101010;
12'b101011100100: data = 6'b101010;
12'b101011100101: data = 6'b101010;
12'b101011100110: data = 6'b101010;
12'b101011100111: data = 6'b101010;
12'b101011101000: data = 6'b101010;
12'b101011101001: data = 6'b101010;
12'b101011101010: data = 6'b101010;
12'b101011101011: data = 6'b101010;
12'b101011101100: data = 6'b101010;
12'b101011101101: data = 6'b101010;
12'b101011101110: data = 6'b101010;
12'b101011101111: data = 6'b101010;
12'b101011110000: data = 6'b101010;
12'b101011110001: data = 6'b101010;
12'b101011110010: data = 6'b101010;
12'b101011110011: data = 6'b101010;
12'b101011110100: data = 6'b101010;
12'b101011110101: data = 6'b101010;
12'b101011110110: data = 6'b101010;
12'b101011110111: data = 6'b101010;
12'b101011111000: data = 6'b101010;
12'b101011111001: data = 6'b101010;
12'b101011111010: data = 6'b101010;
12'b101011111011: data = 6'b101010;
12'b101011111100: data = 6'b101010;
12'b101011111101: data = 6'b101010;
12'b101011111110: data = 6'b101010;
12'b101011111111: data = 6'b101010;
12'b1010111000000: data = 6'b101010;
12'b1010111000001: data = 6'b101010;
12'b1010111000010: data = 6'b101010;
12'b1010111000011: data = 6'b101010;
12'b1010111000100: data = 6'b101010;
12'b1010111000101: data = 6'b101010;
12'b1010111000110: data = 6'b101010;
12'b1010111000111: data = 6'b101010;
12'b1010111001000: data = 6'b101010;
12'b1010111001001: data = 6'b101010;
12'b1010111001010: data = 6'b101010;
12'b1010111001011: data = 6'b101010;
12'b1010111001100: data = 6'b101010;
12'b1010111001101: data = 6'b101010;
12'b1010111001110: data = 6'b101010;
12'b1010111001111: data = 6'b101010;
12'b1010111010000: data = 6'b101010;
12'b1010111010001: data = 6'b101010;
12'b1010111010010: data = 6'b101010;
12'b1010111010011: data = 6'b101010;
12'b1010111010100: data = 6'b101010;
12'b1010111010101: data = 6'b101010;
12'b1010111010110: data = 6'b101010;
12'b1010111010111: data = 6'b101010;
12'b1010111011000: data = 6'b101010;
12'b1010111011001: data = 6'b101010;
12'b1010111011010: data = 6'b101010;
12'b1010111011011: data = 6'b101010;
12'b1010111011100: data = 6'b101010;
12'b1010111011101: data = 6'b101010;
12'b1010111011110: data = 6'b101010;
12'b1010111011111: data = 6'b101010;
12'b1010111100000: data = 6'b101010;
12'b1010111100001: data = 6'b101010;
12'b1010111100010: data = 6'b010101;
12'b1010111100011: data = 6'b101001;
12'b1010111100100: data = 6'b101010;
12'b1010111100101: data = 6'b101010;
12'b1010111100110: data = 6'b101010;
12'b1010111100111: data = 6'b101010;
12'b1010111101000: data = 6'b101010;
12'b1010111101001: data = 6'b101010;
12'b1010111101010: data = 6'b101010;
12'b1010111101011: data = 6'b101010;
12'b1010111101100: data = 6'b101010;
12'b1010111101101: data = 6'b101010;
12'b1010111101110: data = 6'b101010;
12'b1010111101111: data = 6'b101010;
12'b1010111110000: data = 6'b101010;
12'b1010111110001: data = 6'b101010;
12'b1010111110010: data = 6'b101010;
12'b1010111110011: data = 6'b101010;
12'b1010111110100: data = 6'b101010;
12'b1010111110101: data = 6'b101010;
12'b1010111110110: data = 6'b101010;
12'b1010111110111: data = 6'b101010;
12'b1010111111000: data = 6'b101010;
12'b1010111111001: data = 6'b101010;
12'b1010111111010: data = 6'b101010;
12'b1010111111011: data = 6'b101010;
12'b1010111111100: data = 6'b101010;
12'b1010111111101: data = 6'b101010;
12'b1010111111110: data = 6'b101010;
12'b1010111111111: data = 6'b101010;
12'b10101110000000: data = 6'b101010;
12'b10101110000001: data = 6'b101010;
12'b10101110000010: data = 6'b101010;
12'b10101110000011: data = 6'b101010;
12'b10101110000100: data = 6'b101010;
12'b10101110000101: data = 6'b101010;
12'b10101110000110: data = 6'b101010;
12'b10101110000111: data = 6'b101010;
12'b10101110001000: data = 6'b101010;
12'b10101110001001: data = 6'b010101;
12'b10101110001010: data = 6'b010101;
12'b10101110001011: data = 6'b010101;
12'b10101110001100: data = 6'b000000;
12'b10101110001101: data = 6'b000000;
12'b10101110001110: data = 6'b101010;
12'b10101110001111: data = 6'b101010;
12'b10101110010000: data = 6'b101010;
12'b10101110010001: data = 6'b101010;
12'b10101110010010: data = 6'b010101;
12'b10101110010011: data = 6'b010101;
12'b10101110010100: data = 6'b010101;
12'b10101110010101: data = 6'b010101;
12'b10101110010110: data = 6'b010101;
12'b10101110010111: data = 6'b010101;
12'b10101110011000: data = 6'b010101;
12'b10101110011001: data = 6'b010101;
12'b10101110011010: data = 6'b010101;
12'b10101110011011: data = 6'b010101;
12'b10101110011100: data = 6'b010101;
12'b10101110011101: data = 6'b010101;
12'b10101110011110: data = 6'b010101;
12'b10101110011111: data = 6'b010101;
12'b10101110100000: data = 6'b010101;
12'b10101110100001: data = 6'b010101;
12'b10101110100010: data = 6'b010101;
12'b10101110100011: data = 6'b010101;
12'b10101110100100: data = 6'b010101;
12'b10101110100101: data = 6'b010101;
12'b10101110100110: data = 6'b010101;
12'b10101110100111: data = 6'b010101;
12'b10101110101000: data = 6'b010101;
12'b10101110101001: data = 6'b010101;
12'b10101110101010: data = 6'b010101;
12'b101100000000: data = 6'b010101;
12'b101100000001: data = 6'b010101;
12'b101100000010: data = 6'b010101;
12'b101100000011: data = 6'b010101;
12'b101100000100: data = 6'b010101;
12'b101100000101: data = 6'b010101;
12'b101100000110: data = 6'b010101;
12'b101100000111: data = 6'b010101;
12'b101100001000: data = 6'b010101;
12'b101100001001: data = 6'b010101;
12'b101100001010: data = 6'b010101;
12'b101100001011: data = 6'b010101;
12'b101100001100: data = 6'b010101;
12'b101100001101: data = 6'b010101;
12'b101100001110: data = 6'b010101;
12'b101100001111: data = 6'b010101;
12'b101100010000: data = 6'b010101;
12'b101100010001: data = 6'b010101;
12'b101100010010: data = 6'b010101;
12'b101100010011: data = 6'b010101;
12'b101100010100: data = 6'b010101;
12'b101100010101: data = 6'b010101;
12'b101100010110: data = 6'b010101;
12'b101100010111: data = 6'b010101;
12'b101100011000: data = 6'b010101;
12'b101100011001: data = 6'b101010;
12'b101100011010: data = 6'b101010;
12'b101100011011: data = 6'b101010;
12'b101100011100: data = 6'b010101;
12'b101100011101: data = 6'b000000;
12'b101100011110: data = 6'b000000;
12'b101100011111: data = 6'b010101;
12'b101100100000: data = 6'b010101;
12'b101100100001: data = 6'b010101;
12'b101100100010: data = 6'b101010;
12'b101100100011: data = 6'b101010;
12'b101100100100: data = 6'b101010;
12'b101100100101: data = 6'b101010;
12'b101100100110: data = 6'b101010;
12'b101100100111: data = 6'b101010;
12'b101100101000: data = 6'b101010;
12'b101100101001: data = 6'b101010;
12'b101100101010: data = 6'b101010;
12'b101100101011: data = 6'b101010;
12'b101100101100: data = 6'b101010;
12'b101100101101: data = 6'b101010;
12'b101100101110: data = 6'b101010;
12'b101100101111: data = 6'b101010;
12'b101100110000: data = 6'b101010;
12'b101100110001: data = 6'b101010;
12'b101100110010: data = 6'b101010;
12'b101100110011: data = 6'b101010;
12'b101100110100: data = 6'b101010;
12'b101100110101: data = 6'b101010;
12'b101100110110: data = 6'b101010;
12'b101100110111: data = 6'b101010;
12'b101100111000: data = 6'b101010;
12'b101100111001: data = 6'b101010;
12'b101100111010: data = 6'b101010;
12'b101100111011: data = 6'b101010;
12'b101100111100: data = 6'b101010;
12'b101100111101: data = 6'b101010;
12'b101100111110: data = 6'b101010;
12'b101100111111: data = 6'b101010;
12'b1011001000000: data = 6'b101010;
12'b1011001000001: data = 6'b101010;
12'b1011001000010: data = 6'b101010;
12'b1011001000011: data = 6'b101010;
12'b1011001000100: data = 6'b101010;
12'b1011001000101: data = 6'b101010;
12'b1011001000110: data = 6'b101010;
12'b1011001000111: data = 6'b101010;
12'b1011001001000: data = 6'b101010;
12'b1011001001001: data = 6'b101010;
12'b1011001001010: data = 6'b101010;
12'b1011001001011: data = 6'b101010;
12'b1011001001100: data = 6'b101010;
12'b1011001001101: data = 6'b101010;
12'b1011001001110: data = 6'b101010;
12'b1011001001111: data = 6'b101010;
12'b1011001010000: data = 6'b101010;
12'b1011001010001: data = 6'b101010;
12'b1011001010010: data = 6'b101010;
12'b1011001010011: data = 6'b101010;
12'b1011001010100: data = 6'b101010;
12'b1011001010101: data = 6'b101010;
12'b1011001010110: data = 6'b101010;
12'b1011001010111: data = 6'b101010;
12'b1011001011000: data = 6'b101010;
12'b1011001011001: data = 6'b101010;
12'b1011001011010: data = 6'b101010;
12'b1011001011011: data = 6'b101010;
12'b1011001011100: data = 6'b101010;
12'b1011001011101: data = 6'b101010;
12'b1011001011110: data = 6'b101010;
12'b1011001011111: data = 6'b101010;
12'b1011001100000: data = 6'b101010;
12'b1011001100001: data = 6'b101010;
12'b1011001100010: data = 6'b010101;
12'b1011001100011: data = 6'b101001;
12'b1011001100100: data = 6'b101010;
12'b1011001100101: data = 6'b101010;
12'b1011001100110: data = 6'b101010;
12'b1011001100111: data = 6'b101010;
12'b1011001101000: data = 6'b101010;
12'b1011001101001: data = 6'b101010;
12'b1011001101010: data = 6'b101010;
12'b1011001101011: data = 6'b101010;
12'b1011001101100: data = 6'b101010;
12'b1011001101101: data = 6'b101010;
12'b1011001101110: data = 6'b101010;
12'b1011001101111: data = 6'b101010;
12'b1011001110000: data = 6'b101010;
12'b1011001110001: data = 6'b101010;
12'b1011001110010: data = 6'b101010;
12'b1011001110011: data = 6'b101010;
12'b1011001110100: data = 6'b101010;
12'b1011001110101: data = 6'b101010;
12'b1011001110110: data = 6'b101010;
12'b1011001110111: data = 6'b101010;
12'b1011001111000: data = 6'b101010;
12'b1011001111001: data = 6'b101010;
12'b1011001111010: data = 6'b101010;
12'b1011001111011: data = 6'b101010;
12'b1011001111100: data = 6'b101010;
12'b1011001111101: data = 6'b101010;
12'b1011001111110: data = 6'b101010;
12'b1011001111111: data = 6'b101010;
12'b10110010000000: data = 6'b101010;
12'b10110010000001: data = 6'b101010;
12'b10110010000010: data = 6'b101010;
12'b10110010000011: data = 6'b101010;
12'b10110010000100: data = 6'b101010;
12'b10110010000101: data = 6'b101010;
12'b10110010000110: data = 6'b101010;
12'b10110010000111: data = 6'b101010;
12'b10110010001000: data = 6'b101010;
12'b10110010001001: data = 6'b010101;
12'b10110010001010: data = 6'b010101;
12'b10110010001011: data = 6'b010101;
12'b10110010001100: data = 6'b000000;
12'b10110010001101: data = 6'b000000;
12'b10110010001110: data = 6'b101010;
12'b10110010001111: data = 6'b101010;
12'b10110010010000: data = 6'b101010;
12'b10110010010001: data = 6'b101010;
12'b10110010010010: data = 6'b010101;
12'b10110010010011: data = 6'b010101;
12'b10110010010100: data = 6'b010101;
12'b10110010010101: data = 6'b010101;
12'b10110010010110: data = 6'b010101;
12'b10110010010111: data = 6'b010101;
12'b10110010011000: data = 6'b010101;
12'b10110010011001: data = 6'b010101;
12'b10110010011010: data = 6'b010101;
12'b10110010011011: data = 6'b010101;
12'b10110010011100: data = 6'b010101;
12'b10110010011101: data = 6'b010101;
12'b10110010011110: data = 6'b010101;
12'b10110010011111: data = 6'b010101;
12'b10110010100000: data = 6'b010101;
12'b10110010100001: data = 6'b010101;
12'b10110010100010: data = 6'b010101;
12'b10110010100011: data = 6'b010101;
12'b10110010100100: data = 6'b010101;
12'b10110010100101: data = 6'b010101;
12'b10110010100110: data = 6'b010101;
12'b10110010100111: data = 6'b010101;
12'b10110010101000: data = 6'b010101;
12'b10110010101001: data = 6'b010101;
12'b10110010101010: data = 6'b010101;
12'b101101000000: data = 6'b010101;
12'b101101000001: data = 6'b010101;
12'b101101000010: data = 6'b010101;
12'b101101000011: data = 6'b010101;
12'b101101000100: data = 6'b010101;
12'b101101000101: data = 6'b010101;
12'b101101000110: data = 6'b010101;
12'b101101000111: data = 6'b010101;
12'b101101001000: data = 6'b010101;
12'b101101001001: data = 6'b010101;
12'b101101001010: data = 6'b010101;
12'b101101001011: data = 6'b010101;
12'b101101001100: data = 6'b010101;
12'b101101001101: data = 6'b010101;
12'b101101001110: data = 6'b010101;
12'b101101001111: data = 6'b010101;
12'b101101010000: data = 6'b010101;
12'b101101010001: data = 6'b010101;
12'b101101010010: data = 6'b010101;
12'b101101010011: data = 6'b010101;
12'b101101010100: data = 6'b010101;
12'b101101010101: data = 6'b010101;
12'b101101010110: data = 6'b010101;
12'b101101010111: data = 6'b010101;
12'b101101011000: data = 6'b010101;
12'b101101011001: data = 6'b101010;
12'b101101011010: data = 6'b101010;
12'b101101011011: data = 6'b101010;
12'b101101011100: data = 6'b010101;
12'b101101011101: data = 6'b000000;
12'b101101011110: data = 6'b000000;
12'b101101011111: data = 6'b010101;
12'b101101100000: data = 6'b010101;
12'b101101100001: data = 6'b010101;
12'b101101100010: data = 6'b101010;
12'b101101100011: data = 6'b101010;
12'b101101100100: data = 6'b101010;
12'b101101100101: data = 6'b101010;
12'b101101100110: data = 6'b101010;
12'b101101100111: data = 6'b101010;
12'b101101101000: data = 6'b101010;
12'b101101101001: data = 6'b101010;
12'b101101101010: data = 6'b101010;
12'b101101101011: data = 6'b101010;
12'b101101101100: data = 6'b101010;
12'b101101101101: data = 6'b101010;
12'b101101101110: data = 6'b101010;
12'b101101101111: data = 6'b101010;
12'b101101110000: data = 6'b101010;
12'b101101110001: data = 6'b101010;
12'b101101110010: data = 6'b101010;
12'b101101110011: data = 6'b101010;
12'b101101110100: data = 6'b101010;
12'b101101110101: data = 6'b101010;
12'b101101110110: data = 6'b101010;
12'b101101110111: data = 6'b101010;
12'b101101111000: data = 6'b101010;
12'b101101111001: data = 6'b101010;
12'b101101111010: data = 6'b101010;
12'b101101111011: data = 6'b101010;
12'b101101111100: data = 6'b101010;
12'b101101111101: data = 6'b101010;
12'b101101111110: data = 6'b101010;
12'b101101111111: data = 6'b101010;
12'b1011011000000: data = 6'b101010;
12'b1011011000001: data = 6'b101010;
12'b1011011000010: data = 6'b101010;
12'b1011011000011: data = 6'b101010;
12'b1011011000100: data = 6'b101010;
12'b1011011000101: data = 6'b101010;
12'b1011011000110: data = 6'b101010;
12'b1011011000111: data = 6'b101001;
12'b1011011001000: data = 6'b010101;
12'b1011011001001: data = 6'b101010;
12'b1011011001010: data = 6'b101010;
12'b1011011001011: data = 6'b101010;
12'b1011011001100: data = 6'b101010;
12'b1011011001101: data = 6'b101010;
12'b1011011001110: data = 6'b101010;
12'b1011011001111: data = 6'b101010;
12'b1011011010000: data = 6'b101010;
12'b1011011010001: data = 6'b101010;
12'b1011011010010: data = 6'b101010;
12'b1011011010011: data = 6'b101010;
12'b1011011010100: data = 6'b101010;
12'b1011011010101: data = 6'b101010;
12'b1011011010110: data = 6'b101010;
12'b1011011010111: data = 6'b101010;
12'b1011011011000: data = 6'b101010;
12'b1011011011001: data = 6'b101010;
12'b1011011011010: data = 6'b101010;
12'b1011011011011: data = 6'b101010;
12'b1011011011100: data = 6'b101010;
12'b1011011011101: data = 6'b101010;
12'b1011011011110: data = 6'b101010;
12'b1011011011111: data = 6'b101010;
12'b1011011100000: data = 6'b101010;
12'b1011011100001: data = 6'b101010;
12'b1011011100010: data = 6'b010101;
12'b1011011100011: data = 6'b101001;
12'b1011011100100: data = 6'b101010;
12'b1011011100101: data = 6'b101010;
12'b1011011100110: data = 6'b101010;
12'b1011011100111: data = 6'b101010;
12'b1011011101000: data = 6'b101010;
12'b1011011101001: data = 6'b101010;
12'b1011011101010: data = 6'b101010;
12'b1011011101011: data = 6'b101010;
12'b1011011101100: data = 6'b101010;
12'b1011011101101: data = 6'b101010;
12'b1011011101110: data = 6'b101010;
12'b1011011101111: data = 6'b101010;
12'b1011011110000: data = 6'b101010;
12'b1011011110001: data = 6'b101010;
12'b1011011110010: data = 6'b101010;
12'b1011011110011: data = 6'b101010;
12'b1011011110100: data = 6'b101010;
12'b1011011110101: data = 6'b101010;
12'b1011011110110: data = 6'b101010;
12'b1011011110111: data = 6'b101010;
12'b1011011111000: data = 6'b101010;
12'b1011011111001: data = 6'b101010;
12'b1011011111010: data = 6'b101010;
12'b1011011111011: data = 6'b101010;
12'b1011011111100: data = 6'b101010;
12'b1011011111101: data = 6'b101010;
12'b1011011111110: data = 6'b101010;
12'b1011011111111: data = 6'b101010;
12'b10110110000000: data = 6'b101010;
12'b10110110000001: data = 6'b101010;
12'b10110110000010: data = 6'b101010;
12'b10110110000011: data = 6'b101010;
12'b10110110000100: data = 6'b101010;
12'b10110110000101: data = 6'b101010;
12'b10110110000110: data = 6'b101010;
12'b10110110000111: data = 6'b101010;
12'b10110110001000: data = 6'b101010;
12'b10110110001001: data = 6'b010101;
12'b10110110001010: data = 6'b010101;
12'b10110110001011: data = 6'b010101;
12'b10110110001100: data = 6'b000000;
12'b10110110001101: data = 6'b000000;
12'b10110110001110: data = 6'b101010;
12'b10110110001111: data = 6'b101010;
12'b10110110010000: data = 6'b101010;
12'b10110110010001: data = 6'b101010;
12'b10110110010010: data = 6'b010101;
12'b10110110010011: data = 6'b010101;
12'b10110110010100: data = 6'b010101;
12'b10110110010101: data = 6'b010101;
12'b10110110010110: data = 6'b010101;
12'b10110110010111: data = 6'b010101;
12'b10110110011000: data = 6'b010101;
12'b10110110011001: data = 6'b010101;
12'b10110110011010: data = 6'b010101;
12'b10110110011011: data = 6'b010101;
12'b10110110011100: data = 6'b010101;
12'b10110110011101: data = 6'b010101;
12'b10110110011110: data = 6'b010101;
12'b10110110011111: data = 6'b010101;
12'b10110110100000: data = 6'b010101;
12'b10110110100001: data = 6'b010101;
12'b10110110100010: data = 6'b010101;
12'b10110110100011: data = 6'b010101;
12'b10110110100100: data = 6'b010101;
12'b10110110100101: data = 6'b010101;
12'b10110110100110: data = 6'b010101;
12'b10110110100111: data = 6'b010101;
12'b10110110101000: data = 6'b010101;
12'b10110110101001: data = 6'b010101;
12'b10110110101010: data = 6'b010101;
12'b101110000000: data = 6'b010101;
12'b101110000001: data = 6'b010101;
12'b101110000010: data = 6'b010101;
12'b101110000011: data = 6'b010101;
12'b101110000100: data = 6'b010101;
12'b101110000101: data = 6'b010101;
12'b101110000110: data = 6'b010101;
12'b101110000111: data = 6'b010101;
12'b101110001000: data = 6'b010101;
12'b101110001001: data = 6'b010101;
12'b101110001010: data = 6'b010101;
12'b101110001011: data = 6'b010101;
12'b101110001100: data = 6'b010101;
12'b101110001101: data = 6'b010101;
12'b101110001110: data = 6'b010101;
12'b101110001111: data = 6'b010101;
12'b101110010000: data = 6'b010101;
12'b101110010001: data = 6'b010101;
12'b101110010010: data = 6'b010101;
12'b101110010011: data = 6'b010101;
12'b101110010100: data = 6'b010101;
12'b101110010101: data = 6'b010101;
12'b101110010110: data = 6'b010101;
12'b101110010111: data = 6'b010101;
12'b101110011000: data = 6'b010101;
12'b101110011001: data = 6'b101010;
12'b101110011010: data = 6'b101010;
12'b101110011011: data = 6'b101010;
12'b101110011100: data = 6'b010101;
12'b101110011101: data = 6'b000000;
12'b101110011110: data = 6'b000000;
12'b101110011111: data = 6'b010101;
12'b101110100000: data = 6'b010101;
12'b101110100001: data = 6'b010101;
12'b101110100010: data = 6'b101010;
12'b101110100011: data = 6'b101010;
12'b101110100100: data = 6'b101010;
12'b101110100101: data = 6'b101010;
12'b101110100110: data = 6'b101010;
12'b101110100111: data = 6'b101010;
12'b101110101000: data = 6'b101010;
12'b101110101001: data = 6'b101010;
12'b101110101010: data = 6'b101010;
12'b101110101011: data = 6'b101010;
12'b101110101100: data = 6'b101010;
12'b101110101101: data = 6'b101010;
12'b101110101110: data = 6'b101010;
12'b101110101111: data = 6'b101010;
12'b101110110000: data = 6'b101010;
12'b101110110001: data = 6'b101010;
12'b101110110010: data = 6'b101010;
12'b101110110011: data = 6'b101010;
12'b101110110100: data = 6'b101010;
12'b101110110101: data = 6'b101010;
12'b101110110110: data = 6'b101010;
12'b101110110111: data = 6'b101010;
12'b101110111000: data = 6'b101010;
12'b101110111001: data = 6'b101010;
12'b101110111010: data = 6'b101010;
12'b101110111011: data = 6'b101010;
12'b101110111100: data = 6'b101010;
12'b101110111101: data = 6'b101010;
12'b101110111110: data = 6'b101010;
12'b101110111111: data = 6'b101010;
12'b1011101000000: data = 6'b101010;
12'b1011101000001: data = 6'b101010;
12'b1011101000010: data = 6'b101010;
12'b1011101000011: data = 6'b101010;
12'b1011101000100: data = 6'b101010;
12'b1011101000101: data = 6'b101010;
12'b1011101000110: data = 6'b101010;
12'b1011101000111: data = 6'b101001;
12'b1011101001000: data = 6'b010101;
12'b1011101001001: data = 6'b101010;
12'b1011101001010: data = 6'b101010;
12'b1011101001011: data = 6'b101010;
12'b1011101001100: data = 6'b101010;
12'b1011101001101: data = 6'b101010;
12'b1011101001110: data = 6'b101010;
12'b1011101001111: data = 6'b101010;
12'b1011101010000: data = 6'b101010;
12'b1011101010001: data = 6'b101010;
12'b1011101010010: data = 6'b101010;
12'b1011101010011: data = 6'b101010;
12'b1011101010100: data = 6'b101010;
12'b1011101010101: data = 6'b101010;
12'b1011101010110: data = 6'b101010;
12'b1011101010111: data = 6'b101010;
12'b1011101011000: data = 6'b101010;
12'b1011101011001: data = 6'b101010;
12'b1011101011010: data = 6'b101010;
12'b1011101011011: data = 6'b101010;
12'b1011101011100: data = 6'b101010;
12'b1011101011101: data = 6'b101010;
12'b1011101011110: data = 6'b101010;
12'b1011101011111: data = 6'b101010;
12'b1011101100000: data = 6'b101010;
12'b1011101100001: data = 6'b101010;
12'b1011101100010: data = 6'b010101;
12'b1011101100011: data = 6'b101001;
12'b1011101100100: data = 6'b101010;
12'b1011101100101: data = 6'b101010;
12'b1011101100110: data = 6'b101010;
12'b1011101100111: data = 6'b101010;
12'b1011101101000: data = 6'b101010;
12'b1011101101001: data = 6'b101010;
12'b1011101101010: data = 6'b101010;
12'b1011101101011: data = 6'b101010;
12'b1011101101100: data = 6'b101010;
12'b1011101101101: data = 6'b101010;
12'b1011101101110: data = 6'b101010;
12'b1011101101111: data = 6'b101010;
12'b1011101110000: data = 6'b101010;
12'b1011101110001: data = 6'b101010;
12'b1011101110010: data = 6'b101010;
12'b1011101110011: data = 6'b101010;
12'b1011101110100: data = 6'b101010;
12'b1011101110101: data = 6'b101010;
12'b1011101110110: data = 6'b101010;
12'b1011101110111: data = 6'b101010;
12'b1011101111000: data = 6'b101010;
12'b1011101111001: data = 6'b101010;
12'b1011101111010: data = 6'b101010;
12'b1011101111011: data = 6'b101010;
12'b1011101111100: data = 6'b101010;
12'b1011101111101: data = 6'b101010;
12'b1011101111110: data = 6'b101010;
12'b1011101111111: data = 6'b101010;
12'b10111010000000: data = 6'b101010;
12'b10111010000001: data = 6'b101010;
12'b10111010000010: data = 6'b101010;
12'b10111010000011: data = 6'b101010;
12'b10111010000100: data = 6'b101010;
12'b10111010000101: data = 6'b101010;
12'b10111010000110: data = 6'b101010;
12'b10111010000111: data = 6'b101010;
12'b10111010001000: data = 6'b101010;
12'b10111010001001: data = 6'b010101;
12'b10111010001010: data = 6'b010101;
12'b10111010001011: data = 6'b010101;
12'b10111010001100: data = 6'b000000;
12'b10111010001101: data = 6'b000000;
12'b10111010001110: data = 6'b101010;
12'b10111010001111: data = 6'b101010;
12'b10111010010000: data = 6'b101010;
12'b10111010010001: data = 6'b101010;
12'b10111010010010: data = 6'b010101;
12'b10111010010011: data = 6'b010101;
12'b10111010010100: data = 6'b010101;
12'b10111010010101: data = 6'b010101;
12'b10111010010110: data = 6'b010101;
12'b10111010010111: data = 6'b010101;
12'b10111010011000: data = 6'b010101;
12'b10111010011001: data = 6'b010101;
12'b10111010011010: data = 6'b010101;
12'b10111010011011: data = 6'b010101;
12'b10111010011100: data = 6'b010101;
12'b10111010011101: data = 6'b010101;
12'b10111010011110: data = 6'b010101;
12'b10111010011111: data = 6'b010101;
12'b10111010100000: data = 6'b010101;
12'b10111010100001: data = 6'b010101;
12'b10111010100010: data = 6'b010101;
12'b10111010100011: data = 6'b010101;
12'b10111010100100: data = 6'b010101;
12'b10111010100101: data = 6'b010101;
12'b10111010100110: data = 6'b010101;
12'b10111010100111: data = 6'b010101;
12'b10111010101000: data = 6'b010101;
12'b10111010101001: data = 6'b010101;
12'b10111010101010: data = 6'b010101;
12'b101111000000: data = 6'b010101;
12'b101111000001: data = 6'b010101;
12'b101111000010: data = 6'b010101;
12'b101111000011: data = 6'b010101;
12'b101111000100: data = 6'b010101;
12'b101111000101: data = 6'b010101;
12'b101111000110: data = 6'b010101;
12'b101111000111: data = 6'b010101;
12'b101111001000: data = 6'b010101;
12'b101111001001: data = 6'b010101;
12'b101111001010: data = 6'b010101;
12'b101111001011: data = 6'b010101;
12'b101111001100: data = 6'b010101;
12'b101111001101: data = 6'b010101;
12'b101111001110: data = 6'b010101;
12'b101111001111: data = 6'b010101;
12'b101111010000: data = 6'b010101;
12'b101111010001: data = 6'b010101;
12'b101111010010: data = 6'b010101;
12'b101111010011: data = 6'b010101;
12'b101111010100: data = 6'b010101;
12'b101111010101: data = 6'b010101;
12'b101111010110: data = 6'b010101;
12'b101111010111: data = 6'b010101;
12'b101111011000: data = 6'b010101;
12'b101111011001: data = 6'b101010;
12'b101111011010: data = 6'b101010;
12'b101111011011: data = 6'b101010;
12'b101111011100: data = 6'b010101;
12'b101111011101: data = 6'b000000;
12'b101111011110: data = 6'b000000;
12'b101111011111: data = 6'b010101;
12'b101111100000: data = 6'b010101;
12'b101111100001: data = 6'b010101;
12'b101111100010: data = 6'b101010;
12'b101111100011: data = 6'b101010;
12'b101111100100: data = 6'b101010;
12'b101111100101: data = 6'b101010;
12'b101111100110: data = 6'b101010;
12'b101111100111: data = 6'b101010;
12'b101111101000: data = 6'b101010;
12'b101111101001: data = 6'b101010;
12'b101111101010: data = 6'b101010;
12'b101111101011: data = 6'b101010;
12'b101111101100: data = 6'b101010;
12'b101111101101: data = 6'b101010;
12'b101111101110: data = 6'b101010;
12'b101111101111: data = 6'b101010;
12'b101111110000: data = 6'b101010;
12'b101111110001: data = 6'b101010;
12'b101111110010: data = 6'b101010;
12'b101111110011: data = 6'b101010;
12'b101111110100: data = 6'b101010;
12'b101111110101: data = 6'b101010;
12'b101111110110: data = 6'b101010;
12'b101111110111: data = 6'b101010;
12'b101111111000: data = 6'b101010;
12'b101111111001: data = 6'b101010;
12'b101111111010: data = 6'b101010;
12'b101111111011: data = 6'b101010;
12'b101111111100: data = 6'b101010;
12'b101111111101: data = 6'b101010;
12'b101111111110: data = 6'b101010;
12'b101111111111: data = 6'b101010;
12'b1011111000000: data = 6'b101010;
12'b1011111000001: data = 6'b101010;
12'b1011111000010: data = 6'b101010;
12'b1011111000011: data = 6'b101010;
12'b1011111000100: data = 6'b101010;
12'b1011111000101: data = 6'b101010;
12'b1011111000110: data = 6'b101010;
12'b1011111000111: data = 6'b101001;
12'b1011111001000: data = 6'b010101;
12'b1011111001001: data = 6'b101010;
12'b1011111001010: data = 6'b101010;
12'b1011111001011: data = 6'b101010;
12'b1011111001100: data = 6'b101010;
12'b1011111001101: data = 6'b101010;
12'b1011111001110: data = 6'b101010;
12'b1011111001111: data = 6'b101010;
12'b1011111010000: data = 6'b101010;
12'b1011111010001: data = 6'b101010;
12'b1011111010010: data = 6'b101010;
12'b1011111010011: data = 6'b101010;
12'b1011111010100: data = 6'b101010;
12'b1011111010101: data = 6'b101010;
12'b1011111010110: data = 6'b101010;
12'b1011111010111: data = 6'b101010;
12'b1011111011000: data = 6'b101010;
12'b1011111011001: data = 6'b101010;
12'b1011111011010: data = 6'b101010;
12'b1011111011011: data = 6'b101010;
12'b1011111011100: data = 6'b101010;
12'b1011111011101: data = 6'b101010;
12'b1011111011110: data = 6'b101010;
12'b1011111011111: data = 6'b101010;
12'b1011111100000: data = 6'b101010;
12'b1011111100001: data = 6'b101010;
12'b1011111100010: data = 6'b010101;
12'b1011111100011: data = 6'b101001;
12'b1011111100100: data = 6'b101010;
12'b1011111100101: data = 6'b101010;
12'b1011111100110: data = 6'b101010;
12'b1011111100111: data = 6'b101010;
12'b1011111101000: data = 6'b101010;
12'b1011111101001: data = 6'b101010;
12'b1011111101010: data = 6'b101010;
12'b1011111101011: data = 6'b101010;
12'b1011111101100: data = 6'b101010;
12'b1011111101101: data = 6'b101010;
12'b1011111101110: data = 6'b101010;
12'b1011111101111: data = 6'b101010;
12'b1011111110000: data = 6'b101010;
12'b1011111110001: data = 6'b101010;
12'b1011111110010: data = 6'b101010;
12'b1011111110011: data = 6'b101010;
12'b1011111110100: data = 6'b101010;
12'b1011111110101: data = 6'b101010;
12'b1011111110110: data = 6'b101010;
12'b1011111110111: data = 6'b101010;
12'b1011111111000: data = 6'b101010;
12'b1011111111001: data = 6'b101010;
12'b1011111111010: data = 6'b101010;
12'b1011111111011: data = 6'b101010;
12'b1011111111100: data = 6'b101010;
12'b1011111111101: data = 6'b101010;
12'b1011111111110: data = 6'b101010;
12'b1011111111111: data = 6'b101010;
12'b10111110000000: data = 6'b101010;
12'b10111110000001: data = 6'b101010;
12'b10111110000010: data = 6'b101010;
12'b10111110000011: data = 6'b101010;
12'b10111110000100: data = 6'b101010;
12'b10111110000101: data = 6'b101010;
12'b10111110000110: data = 6'b101010;
12'b10111110000111: data = 6'b101010;
12'b10111110001000: data = 6'b101010;
12'b10111110001001: data = 6'b010101;
12'b10111110001010: data = 6'b010101;
12'b10111110001011: data = 6'b010101;
12'b10111110001100: data = 6'b000000;
12'b10111110001101: data = 6'b000000;
12'b10111110001110: data = 6'b101010;
12'b10111110001111: data = 6'b101010;
12'b10111110010000: data = 6'b101010;
12'b10111110010001: data = 6'b101010;
12'b10111110010010: data = 6'b010101;
12'b10111110010011: data = 6'b010101;
12'b10111110010100: data = 6'b010101;
12'b10111110010101: data = 6'b010101;
12'b10111110010110: data = 6'b010101;
12'b10111110010111: data = 6'b010101;
12'b10111110011000: data = 6'b010101;
12'b10111110011001: data = 6'b010101;
12'b10111110011010: data = 6'b010101;
12'b10111110011011: data = 6'b010101;
12'b10111110011100: data = 6'b010101;
12'b10111110011101: data = 6'b010101;
12'b10111110011110: data = 6'b010101;
12'b10111110011111: data = 6'b010101;
12'b10111110100000: data = 6'b010101;
12'b10111110100001: data = 6'b010101;
12'b10111110100010: data = 6'b010101;
12'b10111110100011: data = 6'b010101;
12'b10111110100100: data = 6'b010101;
12'b10111110100101: data = 6'b010101;
12'b10111110100110: data = 6'b010101;
12'b10111110100111: data = 6'b010101;
12'b10111110101000: data = 6'b010101;
12'b10111110101001: data = 6'b010101;
12'b10111110101010: data = 6'b010101;
12'b110000000000: data = 6'b010101;
12'b110000000001: data = 6'b010101;
12'b110000000010: data = 6'b010101;
12'b110000000011: data = 6'b010101;
12'b110000000100: data = 6'b010101;
12'b110000000101: data = 6'b010101;
12'b110000000110: data = 6'b010101;
12'b110000000111: data = 6'b010101;
12'b110000001000: data = 6'b010101;
12'b110000001001: data = 6'b010101;
12'b110000001010: data = 6'b010101;
12'b110000001011: data = 6'b010101;
12'b110000001100: data = 6'b010101;
12'b110000001101: data = 6'b010101;
12'b110000001110: data = 6'b010101;
12'b110000001111: data = 6'b010101;
12'b110000010000: data = 6'b010101;
12'b110000010001: data = 6'b010101;
12'b110000010010: data = 6'b010101;
12'b110000010011: data = 6'b010101;
12'b110000010100: data = 6'b010101;
12'b110000010101: data = 6'b010101;
12'b110000010110: data = 6'b010101;
12'b110000010111: data = 6'b010101;
12'b110000011000: data = 6'b010101;
12'b110000011001: data = 6'b101010;
12'b110000011010: data = 6'b101010;
12'b110000011011: data = 6'b101010;
12'b110000011100: data = 6'b010101;
12'b110000011101: data = 6'b000000;
12'b110000011110: data = 6'b000000;
12'b110000011111: data = 6'b010101;
12'b110000100000: data = 6'b010101;
12'b110000100001: data = 6'b010101;
12'b110000100010: data = 6'b101010;
12'b110000100011: data = 6'b101010;
12'b110000100100: data = 6'b101010;
12'b110000100101: data = 6'b101010;
12'b110000100110: data = 6'b101010;
12'b110000100111: data = 6'b101010;
12'b110000101000: data = 6'b111111;
12'b110000101001: data = 6'b111111;
12'b110000101010: data = 6'b111111;
12'b110000101011: data = 6'b111111;
12'b110000101100: data = 6'b101010;
12'b110000101101: data = 6'b111111;
12'b110000101110: data = 6'b111111;
12'b110000101111: data = 6'b111111;
12'b110000110000: data = 6'b111111;
12'b110000110001: data = 6'b111111;
12'b110000110010: data = 6'b111111;
12'b110000110011: data = 6'b111111;
12'b110000110100: data = 6'b111111;
12'b110000110101: data = 6'b111111;
12'b110000110110: data = 6'b111111;
12'b110000110111: data = 6'b111111;
12'b110000111000: data = 6'b111111;
12'b110000111001: data = 6'b111111;
12'b110000111010: data = 6'b111111;
12'b110000111011: data = 6'b111111;
12'b110000111100: data = 6'b111111;
12'b110000111101: data = 6'b111111;
12'b110000111110: data = 6'b111111;
12'b110000111111: data = 6'b111111;
12'b1100001000000: data = 6'b111111;
12'b1100001000001: data = 6'b101010;
12'b1100001000010: data = 6'b101010;
12'b1100001000011: data = 6'b101010;
12'b1100001000100: data = 6'b101010;
12'b1100001000101: data = 6'b101010;
12'b1100001000110: data = 6'b101010;
12'b1100001000111: data = 6'b101010;
12'b1100001001000: data = 6'b010101;
12'b1100001001001: data = 6'b101010;
12'b1100001001010: data = 6'b111111;
12'b1100001001011: data = 6'b111111;
12'b1100001001100: data = 6'b111111;
12'b1100001001101: data = 6'b111111;
12'b1100001001110: data = 6'b111111;
12'b1100001001111: data = 6'b111111;
12'b1100001010000: data = 6'b111111;
12'b1100001010001: data = 6'b111111;
12'b1100001010010: data = 6'b111111;
12'b1100001010011: data = 6'b111111;
12'b1100001010100: data = 6'b111111;
12'b1100001010101: data = 6'b111111;
12'b1100001010110: data = 6'b111111;
12'b1100001010111: data = 6'b111111;
12'b1100001011000: data = 6'b111111;
12'b1100001011001: data = 6'b111111;
12'b1100001011010: data = 6'b111111;
12'b1100001011011: data = 6'b111111;
12'b1100001011100: data = 6'b111111;
12'b1100001011101: data = 6'b111111;
12'b1100001011110: data = 6'b111111;
12'b1100001011111: data = 6'b111111;
12'b1100001100000: data = 6'b111111;
12'b1100001100001: data = 6'b101010;
12'b1100001100010: data = 6'b010101;
12'b1100001100011: data = 6'b101001;
12'b1100001100100: data = 6'b101010;
12'b1100001100101: data = 6'b101010;
12'b1100001100110: data = 6'b101010;
12'b1100001100111: data = 6'b101010;
12'b1100001101000: data = 6'b101010;
12'b1100001101001: data = 6'b101010;
12'b1100001101010: data = 6'b111111;
12'b1100001101011: data = 6'b111111;
12'b1100001101100: data = 6'b111111;
12'b1100001101101: data = 6'b111111;
12'b1100001101110: data = 6'b111111;
12'b1100001101111: data = 6'b111111;
12'b1100001110000: data = 6'b111111;
12'b1100001110001: data = 6'b111111;
12'b1100001110010: data = 6'b111111;
12'b1100001110011: data = 6'b111111;
12'b1100001110100: data = 6'b111111;
12'b1100001110101: data = 6'b111111;
12'b1100001110110: data = 6'b111111;
12'b1100001110111: data = 6'b111111;
12'b1100001111000: data = 6'b111111;
12'b1100001111001: data = 6'b111111;
12'b1100001111010: data = 6'b111111;
12'b1100001111011: data = 6'b111111;
12'b1100001111100: data = 6'b111111;
12'b1100001111101: data = 6'b111111;
12'b1100001111110: data = 6'b111111;
12'b1100001111111: data = 6'b111111;
12'b11000010000000: data = 6'b111111;
12'b11000010000001: data = 6'b111111;
12'b11000010000010: data = 6'b111111;
12'b11000010000011: data = 6'b101010;
12'b11000010000100: data = 6'b101010;
12'b11000010000101: data = 6'b101010;
12'b11000010000110: data = 6'b101010;
12'b11000010000111: data = 6'b101010;
12'b11000010001000: data = 6'b101010;
12'b11000010001001: data = 6'b010101;
12'b11000010001010: data = 6'b010101;
12'b11000010001011: data = 6'b010101;
12'b11000010001100: data = 6'b000000;
12'b11000010001101: data = 6'b000000;
12'b11000010001110: data = 6'b101010;
12'b11000010001111: data = 6'b101010;
12'b11000010010000: data = 6'b101010;
12'b11000010010001: data = 6'b101010;
12'b11000010010010: data = 6'b010101;
12'b11000010010011: data = 6'b010101;
12'b11000010010100: data = 6'b010101;
12'b11000010010101: data = 6'b010101;
12'b11000010010110: data = 6'b010101;
12'b11000010010111: data = 6'b010101;
12'b11000010011000: data = 6'b010101;
12'b11000010011001: data = 6'b010101;
12'b11000010011010: data = 6'b010101;
12'b11000010011011: data = 6'b010101;
12'b11000010011100: data = 6'b010101;
12'b11000010011101: data = 6'b010101;
12'b11000010011110: data = 6'b010101;
12'b11000010011111: data = 6'b010101;
12'b11000010100000: data = 6'b010101;
12'b11000010100001: data = 6'b010101;
12'b11000010100010: data = 6'b010101;
12'b11000010100011: data = 6'b010101;
12'b11000010100100: data = 6'b010101;
12'b11000010100101: data = 6'b010101;
12'b11000010100110: data = 6'b010101;
12'b11000010100111: data = 6'b010101;
12'b11000010101000: data = 6'b010101;
12'b11000010101001: data = 6'b010101;
12'b11000010101010: data = 6'b010101;
12'b110001000000: data = 6'b010101;
12'b110001000001: data = 6'b010101;
12'b110001000010: data = 6'b010101;
12'b110001000011: data = 6'b010101;
12'b110001000100: data = 6'b010101;
12'b110001000101: data = 6'b010101;
12'b110001000110: data = 6'b010101;
12'b110001000111: data = 6'b010101;
12'b110001001000: data = 6'b010101;
12'b110001001001: data = 6'b010101;
12'b110001001010: data = 6'b010101;
12'b110001001011: data = 6'b010101;
12'b110001001100: data = 6'b010101;
12'b110001001101: data = 6'b010101;
12'b110001001110: data = 6'b010101;
12'b110001001111: data = 6'b010101;
12'b110001010000: data = 6'b010101;
12'b110001010001: data = 6'b010101;
12'b110001010010: data = 6'b010101;
12'b110001010011: data = 6'b010101;
12'b110001010100: data = 6'b010101;
12'b110001010101: data = 6'b010101;
12'b110001010110: data = 6'b010101;
12'b110001010111: data = 6'b010101;
12'b110001011000: data = 6'b010101;
12'b110001011001: data = 6'b101010;
12'b110001011010: data = 6'b101010;
12'b110001011011: data = 6'b101010;
12'b110001011100: data = 6'b010101;
12'b110001011101: data = 6'b000000;
12'b110001011110: data = 6'b000000;
12'b110001011111: data = 6'b010101;
12'b110001100000: data = 6'b010101;
12'b110001100001: data = 6'b010101;
12'b110001100010: data = 6'b101010;
12'b110001100011: data = 6'b101010;
12'b110001100100: data = 6'b101010;
12'b110001100101: data = 6'b101010;
12'b110001100110: data = 6'b101010;
12'b110001100111: data = 6'b101010;
12'b110001101000: data = 6'b111111;
12'b110001101001: data = 6'b111111;
12'b110001101010: data = 6'b111111;
12'b110001101011: data = 6'b111111;
12'b110001101100: data = 6'b111111;
12'b110001101101: data = 6'b111111;
12'b110001101110: data = 6'b111111;
12'b110001101111: data = 6'b111111;
12'b110001110000: data = 6'b111111;
12'b110001110001: data = 6'b111111;
12'b110001110010: data = 6'b111111;
12'b110001110011: data = 6'b111111;
12'b110001110100: data = 6'b111111;
12'b110001110101: data = 6'b111111;
12'b110001110110: data = 6'b111111;
12'b110001110111: data = 6'b111111;
12'b110001111000: data = 6'b111111;
12'b110001111001: data = 6'b111111;
12'b110001111010: data = 6'b111111;
12'b110001111011: data = 6'b111111;
12'b110001111100: data = 6'b111111;
12'b110001111101: data = 6'b111111;
12'b110001111110: data = 6'b111111;
12'b110001111111: data = 6'b111111;
12'b1100011000000: data = 6'b111111;
12'b1100011000001: data = 6'b101010;
12'b1100011000010: data = 6'b101010;
12'b1100011000011: data = 6'b101010;
12'b1100011000100: data = 6'b101010;
12'b1100011000101: data = 6'b101010;
12'b1100011000110: data = 6'b101010;
12'b1100011000111: data = 6'b101010;
12'b1100011001000: data = 6'b101001;
12'b1100011001001: data = 6'b101010;
12'b1100011001010: data = 6'b111111;
12'b1100011001011: data = 6'b111111;
12'b1100011001100: data = 6'b111111;
12'b1100011001101: data = 6'b111111;
12'b1100011001110: data = 6'b111111;
12'b1100011001111: data = 6'b111111;
12'b1100011010000: data = 6'b111111;
12'b1100011010001: data = 6'b111111;
12'b1100011010010: data = 6'b111111;
12'b1100011010011: data = 6'b111111;
12'b1100011010100: data = 6'b111111;
12'b1100011010101: data = 6'b111111;
12'b1100011010110: data = 6'b111111;
12'b1100011010111: data = 6'b111111;
12'b1100011011000: data = 6'b111111;
12'b1100011011001: data = 6'b111111;
12'b1100011011010: data = 6'b111111;
12'b1100011011011: data = 6'b111111;
12'b1100011011100: data = 6'b111111;
12'b1100011011101: data = 6'b111111;
12'b1100011011110: data = 6'b111111;
12'b1100011011111: data = 6'b111111;
12'b1100011100000: data = 6'b111111;
12'b1100011100001: data = 6'b101010;
12'b1100011100010: data = 6'b010101;
12'b1100011100011: data = 6'b101001;
12'b1100011100100: data = 6'b101010;
12'b1100011100101: data = 6'b101010;
12'b1100011100110: data = 6'b101010;
12'b1100011100111: data = 6'b101010;
12'b1100011101000: data = 6'b101010;
12'b1100011101001: data = 6'b101010;
12'b1100011101010: data = 6'b111111;
12'b1100011101011: data = 6'b111111;
12'b1100011101100: data = 6'b111111;
12'b1100011101101: data = 6'b111111;
12'b1100011101110: data = 6'b111111;
12'b1100011101111: data = 6'b111111;
12'b1100011110000: data = 6'b111111;
12'b1100011110001: data = 6'b111111;
12'b1100011110010: data = 6'b111111;
12'b1100011110011: data = 6'b111111;
12'b1100011110100: data = 6'b111111;
12'b1100011110101: data = 6'b111111;
12'b1100011110110: data = 6'b111111;
12'b1100011110111: data = 6'b111111;
12'b1100011111000: data = 6'b111111;
12'b1100011111001: data = 6'b111111;
12'b1100011111010: data = 6'b111111;
12'b1100011111011: data = 6'b111111;
12'b1100011111100: data = 6'b111111;
12'b1100011111101: data = 6'b111111;
12'b1100011111110: data = 6'b111111;
12'b1100011111111: data = 6'b111111;
12'b11000110000000: data = 6'b111111;
12'b11000110000001: data = 6'b111111;
12'b11000110000010: data = 6'b111111;
12'b11000110000011: data = 6'b101010;
12'b11000110000100: data = 6'b101010;
12'b11000110000101: data = 6'b101010;
12'b11000110000110: data = 6'b101010;
12'b11000110000111: data = 6'b101010;
12'b11000110001000: data = 6'b101010;
12'b11000110001001: data = 6'b010101;
12'b11000110001010: data = 6'b010101;
12'b11000110001011: data = 6'b010101;
12'b11000110001100: data = 6'b000000;
12'b11000110001101: data = 6'b000000;
12'b11000110001110: data = 6'b101010;
12'b11000110001111: data = 6'b101010;
12'b11000110010000: data = 6'b101010;
12'b11000110010001: data = 6'b101010;
12'b11000110010010: data = 6'b010101;
12'b11000110010011: data = 6'b010101;
12'b11000110010100: data = 6'b010101;
12'b11000110010101: data = 6'b010101;
12'b11000110010110: data = 6'b010101;
12'b11000110010111: data = 6'b010101;
12'b11000110011000: data = 6'b010101;
12'b11000110011001: data = 6'b010101;
12'b11000110011010: data = 6'b010101;
12'b11000110011011: data = 6'b010101;
12'b11000110011100: data = 6'b010101;
12'b11000110011101: data = 6'b010101;
12'b11000110011110: data = 6'b010101;
12'b11000110011111: data = 6'b010101;
12'b11000110100000: data = 6'b010101;
12'b11000110100001: data = 6'b010101;
12'b11000110100010: data = 6'b010101;
12'b11000110100011: data = 6'b010101;
12'b11000110100100: data = 6'b010101;
12'b11000110100101: data = 6'b010101;
12'b11000110100110: data = 6'b010101;
12'b11000110100111: data = 6'b010101;
12'b11000110101000: data = 6'b010101;
12'b11000110101001: data = 6'b010101;
12'b11000110101010: data = 6'b010101;
12'b110010000000: data = 6'b010101;
12'b110010000001: data = 6'b010101;
12'b110010000010: data = 6'b010101;
12'b110010000011: data = 6'b010101;
12'b110010000100: data = 6'b010101;
12'b110010000101: data = 6'b010101;
12'b110010000110: data = 6'b010101;
12'b110010000111: data = 6'b010101;
12'b110010001000: data = 6'b010101;
12'b110010001001: data = 6'b010101;
12'b110010001010: data = 6'b010101;
12'b110010001011: data = 6'b010101;
12'b110010001100: data = 6'b010101;
12'b110010001101: data = 6'b010101;
12'b110010001110: data = 6'b010101;
12'b110010001111: data = 6'b010101;
12'b110010010000: data = 6'b010101;
12'b110010010001: data = 6'b010101;
12'b110010010010: data = 6'b010101;
12'b110010010011: data = 6'b010101;
12'b110010010100: data = 6'b010101;
12'b110010010101: data = 6'b010101;
12'b110010010110: data = 6'b010101;
12'b110010010111: data = 6'b010101;
12'b110010011000: data = 6'b010101;
12'b110010011001: data = 6'b101010;
12'b110010011010: data = 6'b101010;
12'b110010011011: data = 6'b101010;
12'b110010011100: data = 6'b010101;
12'b110010011101: data = 6'b000000;
12'b110010011110: data = 6'b000000;
12'b110010011111: data = 6'b010101;
12'b110010100000: data = 6'b010101;
12'b110010100001: data = 6'b010101;
12'b110010100010: data = 6'b101010;
12'b110010100011: data = 6'b101010;
12'b110010100100: data = 6'b101010;
12'b110010100101: data = 6'b101010;
12'b110010100110: data = 6'b101010;
12'b110010100111: data = 6'b101010;
12'b110010101000: data = 6'b111111;
12'b110010101001: data = 6'b111111;
12'b110010101010: data = 6'b111111;
12'b110010101011: data = 6'b111111;
12'b110010101100: data = 6'b111111;
12'b110010101101: data = 6'b111111;
12'b110010101110: data = 6'b111111;
12'b110010101111: data = 6'b111111;
12'b110010110000: data = 6'b111111;
12'b110010110001: data = 6'b111111;
12'b110010110010: data = 6'b111111;
12'b110010110011: data = 6'b111111;
12'b110010110100: data = 6'b111111;
12'b110010110101: data = 6'b111111;
12'b110010110110: data = 6'b111111;
12'b110010110111: data = 6'b111111;
12'b110010111000: data = 6'b111111;
12'b110010111001: data = 6'b111111;
12'b110010111010: data = 6'b111111;
12'b110010111011: data = 6'b111111;
12'b110010111100: data = 6'b111111;
12'b110010111101: data = 6'b111111;
12'b110010111110: data = 6'b111111;
12'b110010111111: data = 6'b111111;
12'b1100101000000: data = 6'b111111;
12'b1100101000001: data = 6'b101010;
12'b1100101000010: data = 6'b101010;
12'b1100101000011: data = 6'b101010;
12'b1100101000100: data = 6'b101010;
12'b1100101000101: data = 6'b101010;
12'b1100101000110: data = 6'b101010;
12'b1100101000111: data = 6'b101010;
12'b1100101001000: data = 6'b101010;
12'b1100101001001: data = 6'b101010;
12'b1100101001010: data = 6'b111111;
12'b1100101001011: data = 6'b111111;
12'b1100101001100: data = 6'b111111;
12'b1100101001101: data = 6'b111111;
12'b1100101001110: data = 6'b111111;
12'b1100101001111: data = 6'b111111;
12'b1100101010000: data = 6'b111111;
12'b1100101010001: data = 6'b111111;
12'b1100101010010: data = 6'b111111;
12'b1100101010011: data = 6'b111111;
12'b1100101010100: data = 6'b111111;
12'b1100101010101: data = 6'b111111;
12'b1100101010110: data = 6'b111111;
12'b1100101010111: data = 6'b111111;
12'b1100101011000: data = 6'b111111;
12'b1100101011001: data = 6'b111111;
12'b1100101011010: data = 6'b111111;
12'b1100101011011: data = 6'b111111;
12'b1100101011100: data = 6'b111111;
12'b1100101011101: data = 6'b111111;
12'b1100101011110: data = 6'b111111;
12'b1100101011111: data = 6'b111111;
12'b1100101100000: data = 6'b111111;
12'b1100101100001: data = 6'b101010;
12'b1100101100010: data = 6'b010101;
12'b1100101100011: data = 6'b101010;
12'b1100101100100: data = 6'b101010;
12'b1100101100101: data = 6'b101010;
12'b1100101100110: data = 6'b101010;
12'b1100101100111: data = 6'b101010;
12'b1100101101000: data = 6'b101010;
12'b1100101101001: data = 6'b101010;
12'b1100101101010: data = 6'b111111;
12'b1100101101011: data = 6'b111111;
12'b1100101101100: data = 6'b111111;
12'b1100101101101: data = 6'b111111;
12'b1100101101110: data = 6'b111111;
12'b1100101101111: data = 6'b111111;
12'b1100101110000: data = 6'b111111;
12'b1100101110001: data = 6'b111111;
12'b1100101110010: data = 6'b111111;
12'b1100101110011: data = 6'b111111;
12'b1100101110100: data = 6'b111111;
12'b1100101110101: data = 6'b111111;
12'b1100101110110: data = 6'b111111;
12'b1100101110111: data = 6'b111111;
12'b1100101111000: data = 6'b111111;
12'b1100101111001: data = 6'b111111;
12'b1100101111010: data = 6'b111111;
12'b1100101111011: data = 6'b111111;
12'b1100101111100: data = 6'b111111;
12'b1100101111101: data = 6'b111111;
12'b1100101111110: data = 6'b111111;
12'b1100101111111: data = 6'b111111;
12'b11001010000000: data = 6'b111111;
12'b11001010000001: data = 6'b111111;
12'b11001010000010: data = 6'b111111;
12'b11001010000011: data = 6'b101010;
12'b11001010000100: data = 6'b101010;
12'b11001010000101: data = 6'b101010;
12'b11001010000110: data = 6'b101010;
12'b11001010000111: data = 6'b101010;
12'b11001010001000: data = 6'b101010;
12'b11001010001001: data = 6'b010101;
12'b11001010001010: data = 6'b010101;
12'b11001010001011: data = 6'b010101;
12'b11001010001100: data = 6'b000000;
12'b11001010001101: data = 6'b000000;
12'b11001010001110: data = 6'b101010;
12'b11001010001111: data = 6'b101010;
12'b11001010010000: data = 6'b101010;
12'b11001010010001: data = 6'b101010;
12'b11001010010010: data = 6'b010101;
12'b11001010010011: data = 6'b010101;
12'b11001010010100: data = 6'b010101;
12'b11001010010101: data = 6'b010101;
12'b11001010010110: data = 6'b010101;
12'b11001010010111: data = 6'b010101;
12'b11001010011000: data = 6'b010101;
12'b11001010011001: data = 6'b010101;
12'b11001010011010: data = 6'b010101;
12'b11001010011011: data = 6'b010101;
12'b11001010011100: data = 6'b010101;
12'b11001010011101: data = 6'b010101;
12'b11001010011110: data = 6'b010101;
12'b11001010011111: data = 6'b010101;
12'b11001010100000: data = 6'b010101;
12'b11001010100001: data = 6'b010101;
12'b11001010100010: data = 6'b010101;
12'b11001010100011: data = 6'b010101;
12'b11001010100100: data = 6'b010101;
12'b11001010100101: data = 6'b010101;
12'b11001010100110: data = 6'b010101;
12'b11001010100111: data = 6'b010101;
12'b11001010101000: data = 6'b010101;
12'b11001010101001: data = 6'b010101;
12'b11001010101010: data = 6'b010101;
12'b110011000000: data = 6'b010101;
12'b110011000001: data = 6'b010101;
12'b110011000010: data = 6'b010101;
12'b110011000011: data = 6'b010101;
12'b110011000100: data = 6'b010101;
12'b110011000101: data = 6'b010101;
12'b110011000110: data = 6'b010101;
12'b110011000111: data = 6'b010101;
12'b110011001000: data = 6'b010101;
12'b110011001001: data = 6'b010101;
12'b110011001010: data = 6'b010101;
12'b110011001011: data = 6'b010101;
12'b110011001100: data = 6'b010101;
12'b110011001101: data = 6'b010101;
12'b110011001110: data = 6'b010101;
12'b110011001111: data = 6'b010101;
12'b110011010000: data = 6'b010101;
12'b110011010001: data = 6'b010101;
12'b110011010010: data = 6'b010101;
12'b110011010011: data = 6'b010101;
12'b110011010100: data = 6'b010101;
12'b110011010101: data = 6'b010101;
12'b110011010110: data = 6'b010101;
12'b110011010111: data = 6'b010101;
12'b110011011000: data = 6'b010101;
12'b110011011001: data = 6'b101010;
12'b110011011010: data = 6'b101010;
12'b110011011011: data = 6'b101010;
12'b110011011100: data = 6'b010101;
12'b110011011101: data = 6'b000000;
12'b110011011110: data = 6'b000000;
12'b110011011111: data = 6'b010101;
12'b110011100000: data = 6'b010101;
12'b110011100001: data = 6'b010101;
12'b110011100010: data = 6'b101010;
12'b110011100011: data = 6'b101010;
12'b110011100100: data = 6'b101010;
12'b110011100101: data = 6'b101010;
12'b110011100110: data = 6'b101010;
12'b110011100111: data = 6'b111111;
12'b110011101000: data = 6'b111111;
12'b110011101001: data = 6'b111111;
12'b110011101010: data = 6'b111111;
12'b110011101011: data = 6'b111111;
12'b110011101100: data = 6'b111111;
12'b110011101101: data = 6'b111111;
12'b110011101110: data = 6'b111111;
12'b110011101111: data = 6'b111111;
12'b110011110000: data = 6'b111111;
12'b110011110001: data = 6'b111111;
12'b110011110010: data = 6'b111111;
12'b110011110011: data = 6'b111111;
12'b110011110100: data = 6'b111111;
12'b110011110101: data = 6'b111111;
12'b110011110110: data = 6'b111111;
12'b110011110111: data = 6'b111111;
12'b110011111000: data = 6'b111111;
12'b110011111001: data = 6'b111111;
12'b110011111010: data = 6'b111111;
12'b110011111011: data = 6'b111111;
12'b110011111100: data = 6'b111111;
12'b110011111101: data = 6'b111111;
12'b110011111110: data = 6'b111111;
12'b110011111111: data = 6'b111111;
12'b1100111000000: data = 6'b111111;
12'b1100111000001: data = 6'b111111;
12'b1100111000010: data = 6'b101010;
12'b1100111000011: data = 6'b101010;
12'b1100111000100: data = 6'b101010;
12'b1100111000101: data = 6'b101010;
12'b1100111000110: data = 6'b101010;
12'b1100111000111: data = 6'b101010;
12'b1100111001000: data = 6'b101010;
12'b1100111001001: data = 6'b101010;
12'b1100111001010: data = 6'b111111;
12'b1100111001011: data = 6'b111111;
12'b1100111001100: data = 6'b111111;
12'b1100111001101: data = 6'b111111;
12'b1100111001110: data = 6'b111111;
12'b1100111001111: data = 6'b111111;
12'b1100111010000: data = 6'b111111;
12'b1100111010001: data = 6'b111111;
12'b1100111010010: data = 6'b111111;
12'b1100111010011: data = 6'b111111;
12'b1100111010100: data = 6'b111111;
12'b1100111010101: data = 6'b111111;
12'b1100111010110: data = 6'b111111;
12'b1100111010111: data = 6'b111111;
12'b1100111011000: data = 6'b111111;
12'b1100111011001: data = 6'b111111;
12'b1100111011010: data = 6'b111111;
12'b1100111011011: data = 6'b111111;
12'b1100111011100: data = 6'b111111;
12'b1100111011101: data = 6'b111111;
12'b1100111011110: data = 6'b111111;
12'b1100111011111: data = 6'b111111;
12'b1100111100000: data = 6'b111111;
12'b1100111100001: data = 6'b101010;
12'b1100111100010: data = 6'b101010;
12'b1100111100011: data = 6'b101010;
12'b1100111100100: data = 6'b101010;
12'b1100111100101: data = 6'b101010;
12'b1100111100110: data = 6'b101010;
12'b1100111100111: data = 6'b101010;
12'b1100111101000: data = 6'b101010;
12'b1100111101001: data = 6'b111111;
12'b1100111101010: data = 6'b111111;
12'b1100111101011: data = 6'b111111;
12'b1100111101100: data = 6'b111111;
12'b1100111101101: data = 6'b111111;
12'b1100111101110: data = 6'b111111;
12'b1100111101111: data = 6'b111111;
12'b1100111110000: data = 6'b111111;
12'b1100111110001: data = 6'b111111;
12'b1100111110010: data = 6'b111111;
12'b1100111110011: data = 6'b111111;
12'b1100111110100: data = 6'b111111;
12'b1100111110101: data = 6'b111111;
12'b1100111110110: data = 6'b111111;
12'b1100111110111: data = 6'b111111;
12'b1100111111000: data = 6'b111111;
12'b1100111111001: data = 6'b111111;
12'b1100111111010: data = 6'b111111;
12'b1100111111011: data = 6'b111111;
12'b1100111111100: data = 6'b111111;
12'b1100111111101: data = 6'b111111;
12'b1100111111110: data = 6'b111111;
12'b1100111111111: data = 6'b111111;
12'b11001110000000: data = 6'b111111;
12'b11001110000001: data = 6'b111111;
12'b11001110000010: data = 6'b111111;
12'b11001110000011: data = 6'b111111;
12'b11001110000100: data = 6'b101010;
12'b11001110000101: data = 6'b101010;
12'b11001110000110: data = 6'b101010;
12'b11001110000111: data = 6'b101010;
12'b11001110001000: data = 6'b101010;
12'b11001110001001: data = 6'b010101;
12'b11001110001010: data = 6'b010101;
12'b11001110001011: data = 6'b010101;
12'b11001110001100: data = 6'b000000;
12'b11001110001101: data = 6'b000000;
12'b11001110001110: data = 6'b101010;
12'b11001110001111: data = 6'b101010;
12'b11001110010000: data = 6'b101010;
12'b11001110010001: data = 6'b101010;
12'b11001110010010: data = 6'b010101;
12'b11001110010011: data = 6'b010101;
12'b11001110010100: data = 6'b010101;
12'b11001110010101: data = 6'b010101;
12'b11001110010110: data = 6'b010101;
12'b11001110010111: data = 6'b010101;
12'b11001110011000: data = 6'b010101;
12'b11001110011001: data = 6'b010101;
12'b11001110011010: data = 6'b010101;
12'b11001110011011: data = 6'b010101;
12'b11001110011100: data = 6'b010101;
12'b11001110011101: data = 6'b010101;
12'b11001110011110: data = 6'b010101;
12'b11001110011111: data = 6'b010101;
12'b11001110100000: data = 6'b010101;
12'b11001110100001: data = 6'b010101;
12'b11001110100010: data = 6'b010101;
12'b11001110100011: data = 6'b010101;
12'b11001110100100: data = 6'b010101;
12'b11001110100101: data = 6'b010101;
12'b11001110100110: data = 6'b010101;
12'b11001110100111: data = 6'b010101;
12'b11001110101000: data = 6'b010101;
12'b11001110101001: data = 6'b010101;
12'b11001110101010: data = 6'b010101;
12'b110100000000: data = 6'b010101;
12'b110100000001: data = 6'b010101;
12'b110100000010: data = 6'b010101;
12'b110100000011: data = 6'b010101;
12'b110100000100: data = 6'b010101;
12'b110100000101: data = 6'b010101;
12'b110100000110: data = 6'b010101;
12'b110100000111: data = 6'b010101;
12'b110100001000: data = 6'b010101;
12'b110100001001: data = 6'b010101;
12'b110100001010: data = 6'b010101;
12'b110100001011: data = 6'b010101;
12'b110100001100: data = 6'b010101;
12'b110100001101: data = 6'b010101;
12'b110100001110: data = 6'b010101;
12'b110100001111: data = 6'b010101;
12'b110100010000: data = 6'b010101;
12'b110100010001: data = 6'b010101;
12'b110100010010: data = 6'b010101;
12'b110100010011: data = 6'b010101;
12'b110100010100: data = 6'b010101;
12'b110100010101: data = 6'b010101;
12'b110100010110: data = 6'b010101;
12'b110100010111: data = 6'b010101;
12'b110100011000: data = 6'b010101;
12'b110100011001: data = 6'b101010;
12'b110100011010: data = 6'b101010;
12'b110100011011: data = 6'b101010;
12'b110100011100: data = 6'b010101;
12'b110100011101: data = 6'b000000;
12'b110100011110: data = 6'b000000;
12'b110100011111: data = 6'b010101;
12'b110100100000: data = 6'b010101;
12'b110100100001: data = 6'b010101;
12'b110100100010: data = 6'b101010;
12'b110100100011: data = 6'b101010;
12'b110100100100: data = 6'b101010;
12'b110100100101: data = 6'b101010;
12'b110100100110: data = 6'b101010;
12'b110100100111: data = 6'b111111;
12'b110100101000: data = 6'b111111;
12'b110100101001: data = 6'b111111;
12'b110100101010: data = 6'b111111;
12'b110100101011: data = 6'b111111;
12'b110100101100: data = 6'b111111;
12'b110100101101: data = 6'b111111;
12'b110100101110: data = 6'b111111;
12'b110100101111: data = 6'b111111;
12'b110100110000: data = 6'b111111;
12'b110100110001: data = 6'b111111;
12'b110100110010: data = 6'b111111;
12'b110100110011: data = 6'b111111;
12'b110100110100: data = 6'b111111;
12'b110100110101: data = 6'b111111;
12'b110100110110: data = 6'b111111;
12'b110100110111: data = 6'b111111;
12'b110100111000: data = 6'b111111;
12'b110100111001: data = 6'b111111;
12'b110100111010: data = 6'b111111;
12'b110100111011: data = 6'b111111;
12'b110100111100: data = 6'b111111;
12'b110100111101: data = 6'b111111;
12'b110100111110: data = 6'b111111;
12'b110100111111: data = 6'b111111;
12'b1101001000000: data = 6'b111111;
12'b1101001000001: data = 6'b111111;
12'b1101001000010: data = 6'b101010;
12'b1101001000011: data = 6'b101010;
12'b1101001000100: data = 6'b101010;
12'b1101001000101: data = 6'b101010;
12'b1101001000110: data = 6'b101010;
12'b1101001000111: data = 6'b101010;
12'b1101001001000: data = 6'b101010;
12'b1101001001001: data = 6'b101010;
12'b1101001001010: data = 6'b111111;
12'b1101001001011: data = 6'b111111;
12'b1101001001100: data = 6'b111111;
12'b1101001001101: data = 6'b111111;
12'b1101001001110: data = 6'b111111;
12'b1101001001111: data = 6'b111111;
12'b1101001010000: data = 6'b111111;
12'b1101001010001: data = 6'b111111;
12'b1101001010010: data = 6'b111111;
12'b1101001010011: data = 6'b111111;
12'b1101001010100: data = 6'b111111;
12'b1101001010101: data = 6'b111111;
12'b1101001010110: data = 6'b111111;
12'b1101001010111: data = 6'b111111;
12'b1101001011000: data = 6'b111111;
12'b1101001011001: data = 6'b111111;
12'b1101001011010: data = 6'b111111;
12'b1101001011011: data = 6'b111111;
12'b1101001011100: data = 6'b111111;
12'b1101001011101: data = 6'b111111;
12'b1101001011110: data = 6'b111111;
12'b1101001011111: data = 6'b111111;
12'b1101001100000: data = 6'b111111;
12'b1101001100001: data = 6'b101010;
12'b1101001100010: data = 6'b101010;
12'b1101001100011: data = 6'b101010;
12'b1101001100100: data = 6'b101010;
12'b1101001100101: data = 6'b101010;
12'b1101001100110: data = 6'b101010;
12'b1101001100111: data = 6'b101010;
12'b1101001101000: data = 6'b101010;
12'b1101001101001: data = 6'b111111;
12'b1101001101010: data = 6'b111111;
12'b1101001101011: data = 6'b111111;
12'b1101001101100: data = 6'b111111;
12'b1101001101101: data = 6'b111111;
12'b1101001101110: data = 6'b111111;
12'b1101001101111: data = 6'b111111;
12'b1101001110000: data = 6'b111111;
12'b1101001110001: data = 6'b111111;
12'b1101001110010: data = 6'b111111;
12'b1101001110011: data = 6'b111111;
12'b1101001110100: data = 6'b111111;
12'b1101001110101: data = 6'b111111;
12'b1101001110110: data = 6'b111111;
12'b1101001110111: data = 6'b111111;
12'b1101001111000: data = 6'b111111;
12'b1101001111001: data = 6'b111111;
12'b1101001111010: data = 6'b111111;
12'b1101001111011: data = 6'b111111;
12'b1101001111100: data = 6'b111111;
12'b1101001111101: data = 6'b111111;
12'b1101001111110: data = 6'b111111;
12'b1101001111111: data = 6'b111111;
12'b11010010000000: data = 6'b111111;
12'b11010010000001: data = 6'b111111;
12'b11010010000010: data = 6'b111111;
12'b11010010000011: data = 6'b111111;
12'b11010010000100: data = 6'b101010;
12'b11010010000101: data = 6'b101010;
12'b11010010000110: data = 6'b101010;
12'b11010010000111: data = 6'b101010;
12'b11010010001000: data = 6'b101010;
12'b11010010001001: data = 6'b010101;
12'b11010010001010: data = 6'b010101;
12'b11010010001011: data = 6'b010101;
12'b11010010001100: data = 6'b000000;
12'b11010010001101: data = 6'b000000;
12'b11010010001110: data = 6'b101010;
12'b11010010001111: data = 6'b101010;
12'b11010010010000: data = 6'b101010;
12'b11010010010001: data = 6'b101010;
12'b11010010010010: data = 6'b010101;
12'b11010010010011: data = 6'b010101;
12'b11010010010100: data = 6'b010101;
12'b11010010010101: data = 6'b010101;
12'b11010010010110: data = 6'b010101;
12'b11010010010111: data = 6'b010101;
12'b11010010011000: data = 6'b010101;
12'b11010010011001: data = 6'b010101;
12'b11010010011010: data = 6'b010101;
12'b11010010011011: data = 6'b010101;
12'b11010010011100: data = 6'b010101;
12'b11010010011101: data = 6'b010101;
12'b11010010011110: data = 6'b010101;
12'b11010010011111: data = 6'b010101;
12'b11010010100000: data = 6'b010101;
12'b11010010100001: data = 6'b010101;
12'b11010010100010: data = 6'b010101;
12'b11010010100011: data = 6'b010101;
12'b11010010100100: data = 6'b010101;
12'b11010010100101: data = 6'b010101;
12'b11010010100110: data = 6'b010101;
12'b11010010100111: data = 6'b010101;
12'b11010010101000: data = 6'b010101;
12'b11010010101001: data = 6'b010101;
12'b11010010101010: data = 6'b010101;
12'b110101000000: data = 6'b010101;
12'b110101000001: data = 6'b010101;
12'b110101000010: data = 6'b010101;
12'b110101000011: data = 6'b010101;
12'b110101000100: data = 6'b010101;
12'b110101000101: data = 6'b010101;
12'b110101000110: data = 6'b010101;
12'b110101000111: data = 6'b010101;
12'b110101001000: data = 6'b010101;
12'b110101001001: data = 6'b010101;
12'b110101001010: data = 6'b010101;
12'b110101001011: data = 6'b010101;
12'b110101001100: data = 6'b010101;
12'b110101001101: data = 6'b010101;
12'b110101001110: data = 6'b010101;
12'b110101001111: data = 6'b010101;
12'b110101010000: data = 6'b010101;
12'b110101010001: data = 6'b010101;
12'b110101010010: data = 6'b010101;
12'b110101010011: data = 6'b010101;
12'b110101010100: data = 6'b010101;
12'b110101010101: data = 6'b010101;
12'b110101010110: data = 6'b010101;
12'b110101010111: data = 6'b010101;
12'b110101011000: data = 6'b010101;
12'b110101011001: data = 6'b101010;
12'b110101011010: data = 6'b101010;
12'b110101011011: data = 6'b101010;
12'b110101011100: data = 6'b010101;
12'b110101011101: data = 6'b000000;
12'b110101011110: data = 6'b000000;
12'b110101011111: data = 6'b010101;
12'b110101100000: data = 6'b010101;
12'b110101100001: data = 6'b010101;
12'b110101100010: data = 6'b101010;
12'b110101100011: data = 6'b101010;
12'b110101100100: data = 6'b101010;
12'b110101100101: data = 6'b101010;
12'b110101100110: data = 6'b101010;
12'b110101100111: data = 6'b111111;
12'b110101101000: data = 6'b111111;
12'b110101101001: data = 6'b111111;
12'b110101101010: data = 6'b111111;
12'b110101101011: data = 6'b111111;
12'b110101101100: data = 6'b111111;
12'b110101101101: data = 6'b111111;
12'b110101101110: data = 6'b111111;
12'b110101101111: data = 6'b111111;
12'b110101110000: data = 6'b111111;
12'b110101110001: data = 6'b111111;
12'b110101110010: data = 6'b111111;
12'b110101110011: data = 6'b111111;
12'b110101110100: data = 6'b111111;
12'b110101110101: data = 6'b111111;
12'b110101110110: data = 6'b111111;
12'b110101110111: data = 6'b111111;
12'b110101111000: data = 6'b111111;
12'b110101111001: data = 6'b111111;
12'b110101111010: data = 6'b111111;
12'b110101111011: data = 6'b111111;
12'b110101111100: data = 6'b111111;
12'b110101111101: data = 6'b111111;
12'b110101111110: data = 6'b111111;
12'b110101111111: data = 6'b111111;
12'b1101011000000: data = 6'b111111;
12'b1101011000001: data = 6'b111111;
12'b1101011000010: data = 6'b101010;
12'b1101011000011: data = 6'b101010;
12'b1101011000100: data = 6'b101010;
12'b1101011000101: data = 6'b101010;
12'b1101011000110: data = 6'b101010;
12'b1101011000111: data = 6'b101010;
12'b1101011001000: data = 6'b101010;
12'b1101011001001: data = 6'b101010;
12'b1101011001010: data = 6'b111111;
12'b1101011001011: data = 6'b111111;
12'b1101011001100: data = 6'b111111;
12'b1101011001101: data = 6'b111111;
12'b1101011001110: data = 6'b111111;
12'b1101011001111: data = 6'b111111;
12'b1101011010000: data = 6'b111111;
12'b1101011010001: data = 6'b111111;
12'b1101011010010: data = 6'b111111;
12'b1101011010011: data = 6'b111111;
12'b1101011010100: data = 6'b111111;
12'b1101011010101: data = 6'b111111;
12'b1101011010110: data = 6'b111111;
12'b1101011010111: data = 6'b111111;
12'b1101011011000: data = 6'b111111;
12'b1101011011001: data = 6'b111111;
12'b1101011011010: data = 6'b111111;
12'b1101011011011: data = 6'b111111;
12'b1101011011100: data = 6'b111111;
12'b1101011011101: data = 6'b111111;
12'b1101011011110: data = 6'b111111;
12'b1101011011111: data = 6'b111111;
12'b1101011100000: data = 6'b111111;
12'b1101011100001: data = 6'b101010;
12'b1101011100010: data = 6'b101010;
12'b1101011100011: data = 6'b101010;
12'b1101011100100: data = 6'b101010;
12'b1101011100101: data = 6'b101010;
12'b1101011100110: data = 6'b101010;
12'b1101011100111: data = 6'b101010;
12'b1101011101000: data = 6'b101010;
12'b1101011101001: data = 6'b111111;
12'b1101011101010: data = 6'b111111;
12'b1101011101011: data = 6'b111111;
12'b1101011101100: data = 6'b111111;
12'b1101011101101: data = 6'b111111;
12'b1101011101110: data = 6'b111111;
12'b1101011101111: data = 6'b111111;
12'b1101011110000: data = 6'b111111;
12'b1101011110001: data = 6'b111111;
12'b1101011110010: data = 6'b111111;
12'b1101011110011: data = 6'b111111;
12'b1101011110100: data = 6'b111111;
12'b1101011110101: data = 6'b111111;
12'b1101011110110: data = 6'b111111;
12'b1101011110111: data = 6'b111111;
12'b1101011111000: data = 6'b111111;
12'b1101011111001: data = 6'b111111;
12'b1101011111010: data = 6'b111111;
12'b1101011111011: data = 6'b111111;
12'b1101011111100: data = 6'b111111;
12'b1101011111101: data = 6'b111111;
12'b1101011111110: data = 6'b111111;
12'b1101011111111: data = 6'b111111;
12'b11010110000000: data = 6'b111111;
12'b11010110000001: data = 6'b111111;
12'b11010110000010: data = 6'b111111;
12'b11010110000011: data = 6'b111111;
12'b11010110000100: data = 6'b101010;
12'b11010110000101: data = 6'b101010;
12'b11010110000110: data = 6'b101010;
12'b11010110000111: data = 6'b101010;
12'b11010110001000: data = 6'b101010;
12'b11010110001001: data = 6'b010101;
12'b11010110001010: data = 6'b010101;
12'b11010110001011: data = 6'b010101;
12'b11010110001100: data = 6'b000000;
12'b11010110001101: data = 6'b000000;
12'b11010110001110: data = 6'b101010;
12'b11010110001111: data = 6'b101010;
12'b11010110010000: data = 6'b101010;
12'b11010110010001: data = 6'b101010;
12'b11010110010010: data = 6'b010101;
12'b11010110010011: data = 6'b010101;
12'b11010110010100: data = 6'b010101;
12'b11010110010101: data = 6'b010101;
12'b11010110010110: data = 6'b010101;
12'b11010110010111: data = 6'b010101;
12'b11010110011000: data = 6'b010101;
12'b11010110011001: data = 6'b010101;
12'b11010110011010: data = 6'b010101;
12'b11010110011011: data = 6'b010101;
12'b11010110011100: data = 6'b010101;
12'b11010110011101: data = 6'b010101;
12'b11010110011110: data = 6'b010101;
12'b11010110011111: data = 6'b010101;
12'b11010110100000: data = 6'b010101;
12'b11010110100001: data = 6'b010101;
12'b11010110100010: data = 6'b010101;
12'b11010110100011: data = 6'b010101;
12'b11010110100100: data = 6'b010101;
12'b11010110100101: data = 6'b010101;
12'b11010110100110: data = 6'b010101;
12'b11010110100111: data = 6'b010101;
12'b11010110101000: data = 6'b010101;
12'b11010110101001: data = 6'b010101;
12'b11010110101010: data = 6'b010101;
12'b110110000000: data = 6'b010101;
12'b110110000001: data = 6'b010101;
12'b110110000010: data = 6'b010101;
12'b110110000011: data = 6'b010101;
12'b110110000100: data = 6'b010101;
12'b110110000101: data = 6'b010101;
12'b110110000110: data = 6'b010101;
12'b110110000111: data = 6'b010101;
12'b110110001000: data = 6'b010101;
12'b110110001001: data = 6'b010101;
12'b110110001010: data = 6'b010101;
12'b110110001011: data = 6'b010101;
12'b110110001100: data = 6'b010101;
12'b110110001101: data = 6'b010101;
12'b110110001110: data = 6'b010101;
12'b110110001111: data = 6'b010101;
12'b110110010000: data = 6'b010101;
12'b110110010001: data = 6'b010101;
12'b110110010010: data = 6'b010101;
12'b110110010011: data = 6'b010101;
12'b110110010100: data = 6'b010101;
12'b110110010101: data = 6'b010101;
12'b110110010110: data = 6'b010101;
12'b110110010111: data = 6'b010101;
12'b110110011000: data = 6'b010101;
12'b110110011001: data = 6'b101010;
12'b110110011010: data = 6'b101010;
12'b110110011011: data = 6'b101010;
12'b110110011100: data = 6'b010101;
12'b110110011101: data = 6'b000000;
12'b110110011110: data = 6'b000000;
12'b110110011111: data = 6'b010101;
12'b110110100000: data = 6'b010101;
12'b110110100001: data = 6'b010101;
12'b110110100010: data = 6'b101010;
12'b110110100011: data = 6'b101010;
12'b110110100100: data = 6'b101010;
12'b110110100101: data = 6'b101010;
12'b110110100110: data = 6'b101010;
12'b110110100111: data = 6'b111111;
12'b110110101000: data = 6'b111111;
12'b110110101001: data = 6'b111111;
12'b110110101010: data = 6'b111111;
12'b110110101011: data = 6'b111111;
12'b110110101100: data = 6'b111111;
12'b110110101101: data = 6'b111111;
12'b110110101110: data = 6'b111111;
12'b110110101111: data = 6'b111111;
12'b110110110000: data = 6'b111111;
12'b110110110001: data = 6'b111111;
12'b110110110010: data = 6'b111111;
12'b110110110011: data = 6'b111111;
12'b110110110100: data = 6'b111111;
12'b110110110101: data = 6'b111111;
12'b110110110110: data = 6'b111111;
12'b110110110111: data = 6'b111111;
12'b110110111000: data = 6'b111111;
12'b110110111001: data = 6'b111111;
12'b110110111010: data = 6'b111111;
12'b110110111011: data = 6'b111111;
12'b110110111100: data = 6'b111111;
12'b110110111101: data = 6'b111111;
12'b110110111110: data = 6'b111111;
12'b110110111111: data = 6'b111111;
12'b1101101000000: data = 6'b111111;
12'b1101101000001: data = 6'b111111;
12'b1101101000010: data = 6'b101010;
12'b1101101000011: data = 6'b101010;
12'b1101101000100: data = 6'b101010;
12'b1101101000101: data = 6'b101010;
12'b1101101000110: data = 6'b101010;
12'b1101101000111: data = 6'b101010;
12'b1101101001000: data = 6'b101010;
12'b1101101001001: data = 6'b101010;
12'b1101101001010: data = 6'b111111;
12'b1101101001011: data = 6'b111111;
12'b1101101001100: data = 6'b111111;
12'b1101101001101: data = 6'b111111;
12'b1101101001110: data = 6'b111111;
12'b1101101001111: data = 6'b111111;
12'b1101101010000: data = 6'b111111;
12'b1101101010001: data = 6'b111111;
12'b1101101010010: data = 6'b111111;
12'b1101101010011: data = 6'b111111;
12'b1101101010100: data = 6'b111111;
12'b1101101010101: data = 6'b111111;
12'b1101101010110: data = 6'b111111;
12'b1101101010111: data = 6'b111111;
12'b1101101011000: data = 6'b111111;
12'b1101101011001: data = 6'b111111;
12'b1101101011010: data = 6'b111111;
12'b1101101011011: data = 6'b111111;
12'b1101101011100: data = 6'b111111;
12'b1101101011101: data = 6'b111111;
12'b1101101011110: data = 6'b111111;
12'b1101101011111: data = 6'b111111;
12'b1101101100000: data = 6'b111111;
12'b1101101100001: data = 6'b101010;
12'b1101101100010: data = 6'b101010;
12'b1101101100011: data = 6'b101010;
12'b1101101100100: data = 6'b101010;
12'b1101101100101: data = 6'b101010;
12'b1101101100110: data = 6'b101010;
12'b1101101100111: data = 6'b101010;
12'b1101101101000: data = 6'b101010;
12'b1101101101001: data = 6'b111111;
12'b1101101101010: data = 6'b111111;
12'b1101101101011: data = 6'b111111;
12'b1101101101100: data = 6'b111111;
12'b1101101101101: data = 6'b111111;
12'b1101101101110: data = 6'b111111;
12'b1101101101111: data = 6'b111111;
12'b1101101110000: data = 6'b111111;
12'b1101101110001: data = 6'b111111;
12'b1101101110010: data = 6'b111111;
12'b1101101110011: data = 6'b111111;
12'b1101101110100: data = 6'b111111;
12'b1101101110101: data = 6'b111111;
12'b1101101110110: data = 6'b111111;
12'b1101101110111: data = 6'b111111;
12'b1101101111000: data = 6'b111111;
12'b1101101111001: data = 6'b111111;
12'b1101101111010: data = 6'b111111;
12'b1101101111011: data = 6'b111111;
12'b1101101111100: data = 6'b111111;
12'b1101101111101: data = 6'b111111;
12'b1101101111110: data = 6'b111111;
12'b1101101111111: data = 6'b111111;
12'b11011010000000: data = 6'b111111;
12'b11011010000001: data = 6'b111111;
12'b11011010000010: data = 6'b111111;
12'b11011010000011: data = 6'b111111;
12'b11011010000100: data = 6'b101010;
12'b11011010000101: data = 6'b101010;
12'b11011010000110: data = 6'b101010;
12'b11011010000111: data = 6'b101010;
12'b11011010001000: data = 6'b101010;
12'b11011010001001: data = 6'b010101;
12'b11011010001010: data = 6'b010101;
12'b11011010001011: data = 6'b010101;
12'b11011010001100: data = 6'b000000;
12'b11011010001101: data = 6'b000000;
12'b11011010001110: data = 6'b101010;
12'b11011010001111: data = 6'b101010;
12'b11011010010000: data = 6'b101010;
12'b11011010010001: data = 6'b101010;
12'b11011010010010: data = 6'b010101;
12'b11011010010011: data = 6'b010101;
12'b11011010010100: data = 6'b010101;
12'b11011010010101: data = 6'b010101;
12'b11011010010110: data = 6'b010101;
12'b11011010010111: data = 6'b010101;
12'b11011010011000: data = 6'b010101;
12'b11011010011001: data = 6'b010101;
12'b11011010011010: data = 6'b010101;
12'b11011010011011: data = 6'b010101;
12'b11011010011100: data = 6'b010101;
12'b11011010011101: data = 6'b010101;
12'b11011010011110: data = 6'b010101;
12'b11011010011111: data = 6'b010101;
12'b11011010100000: data = 6'b010101;
12'b11011010100001: data = 6'b010101;
12'b11011010100010: data = 6'b010101;
12'b11011010100011: data = 6'b010101;
12'b11011010100100: data = 6'b010101;
12'b11011010100101: data = 6'b010101;
12'b11011010100110: data = 6'b010101;
12'b11011010100111: data = 6'b010101;
12'b11011010101000: data = 6'b010101;
12'b11011010101001: data = 6'b010101;
12'b11011010101010: data = 6'b010101;
12'b110111000000: data = 6'b010101;
12'b110111000001: data = 6'b010101;
12'b110111000010: data = 6'b010101;
12'b110111000011: data = 6'b010101;
12'b110111000100: data = 6'b010101;
12'b110111000101: data = 6'b010101;
12'b110111000110: data = 6'b010101;
12'b110111000111: data = 6'b010101;
12'b110111001000: data = 6'b010101;
12'b110111001001: data = 6'b010101;
12'b110111001010: data = 6'b010101;
12'b110111001011: data = 6'b010101;
12'b110111001100: data = 6'b010101;
12'b110111001101: data = 6'b010101;
12'b110111001110: data = 6'b010101;
12'b110111001111: data = 6'b010101;
12'b110111010000: data = 6'b010101;
12'b110111010001: data = 6'b010101;
12'b110111010010: data = 6'b010101;
12'b110111010011: data = 6'b010101;
12'b110111010100: data = 6'b010101;
12'b110111010101: data = 6'b010101;
12'b110111010110: data = 6'b010101;
12'b110111010111: data = 6'b010101;
12'b110111011000: data = 6'b010101;
12'b110111011001: data = 6'b101010;
12'b110111011010: data = 6'b101010;
12'b110111011011: data = 6'b101010;
12'b110111011100: data = 6'b010101;
12'b110111011101: data = 6'b000000;
12'b110111011110: data = 6'b000000;
12'b110111011111: data = 6'b010101;
12'b110111100000: data = 6'b010101;
12'b110111100001: data = 6'b010101;
12'b110111100010: data = 6'b101010;
12'b110111100011: data = 6'b101010;
12'b110111100100: data = 6'b101010;
12'b110111100101: data = 6'b101010;
12'b110111100110: data = 6'b101010;
12'b110111100111: data = 6'b111111;
12'b110111101000: data = 6'b111111;
12'b110111101001: data = 6'b111111;
12'b110111101010: data = 6'b111111;
12'b110111101011: data = 6'b111111;
12'b110111101100: data = 6'b111111;
12'b110111101101: data = 6'b111111;
12'b110111101110: data = 6'b111111;
12'b110111101111: data = 6'b111111;
12'b110111110000: data = 6'b111111;
12'b110111110001: data = 6'b111111;
12'b110111110010: data = 6'b111111;
12'b110111110011: data = 6'b111111;
12'b110111110100: data = 6'b111111;
12'b110111110101: data = 6'b111111;
12'b110111110110: data = 6'b111111;
12'b110111110111: data = 6'b111111;
12'b110111111000: data = 6'b111111;
12'b110111111001: data = 6'b111111;
12'b110111111010: data = 6'b111111;
12'b110111111011: data = 6'b111111;
12'b110111111100: data = 6'b111111;
12'b110111111101: data = 6'b111111;
12'b110111111110: data = 6'b111111;
12'b110111111111: data = 6'b111111;
12'b1101111000000: data = 6'b111111;
12'b1101111000001: data = 6'b111111;
12'b1101111000010: data = 6'b101010;
12'b1101111000011: data = 6'b101010;
12'b1101111000100: data = 6'b101010;
12'b1101111000101: data = 6'b101010;
12'b1101111000110: data = 6'b101010;
12'b1101111000111: data = 6'b101010;
12'b1101111001000: data = 6'b101010;
12'b1101111001001: data = 6'b101010;
12'b1101111001010: data = 6'b111111;
12'b1101111001011: data = 6'b111111;
12'b1101111001100: data = 6'b111111;
12'b1101111001101: data = 6'b111111;
12'b1101111001110: data = 6'b111111;
12'b1101111001111: data = 6'b111111;
12'b1101111010000: data = 6'b111111;
12'b1101111010001: data = 6'b111111;
12'b1101111010010: data = 6'b111111;
12'b1101111010011: data = 6'b111111;
12'b1101111010100: data = 6'b111111;
12'b1101111010101: data = 6'b111111;
12'b1101111010110: data = 6'b111111;
12'b1101111010111: data = 6'b111111;
12'b1101111011000: data = 6'b111111;
12'b1101111011001: data = 6'b111111;
12'b1101111011010: data = 6'b111111;
12'b1101111011011: data = 6'b111111;
12'b1101111011100: data = 6'b111111;
12'b1101111011101: data = 6'b111111;
12'b1101111011110: data = 6'b111111;
12'b1101111011111: data = 6'b111111;
12'b1101111100000: data = 6'b111111;
12'b1101111100001: data = 6'b101010;
12'b1101111100010: data = 6'b101010;
12'b1101111100011: data = 6'b101010;
12'b1101111100100: data = 6'b101010;
12'b1101111100101: data = 6'b101010;
12'b1101111100110: data = 6'b101010;
12'b1101111100111: data = 6'b101010;
12'b1101111101000: data = 6'b101010;
12'b1101111101001: data = 6'b111111;
12'b1101111101010: data = 6'b111111;
12'b1101111101011: data = 6'b111111;
12'b1101111101100: data = 6'b111111;
12'b1101111101101: data = 6'b111111;
12'b1101111101110: data = 6'b111111;
12'b1101111101111: data = 6'b111111;
12'b1101111110000: data = 6'b111111;
12'b1101111110001: data = 6'b111111;
12'b1101111110010: data = 6'b111111;
12'b1101111110011: data = 6'b111111;
12'b1101111110100: data = 6'b111111;
12'b1101111110101: data = 6'b111111;
12'b1101111110110: data = 6'b111111;
12'b1101111110111: data = 6'b111111;
12'b1101111111000: data = 6'b111111;
12'b1101111111001: data = 6'b111111;
12'b1101111111010: data = 6'b111111;
12'b1101111111011: data = 6'b111111;
12'b1101111111100: data = 6'b111111;
12'b1101111111101: data = 6'b111111;
12'b1101111111110: data = 6'b111111;
12'b1101111111111: data = 6'b111111;
12'b11011110000000: data = 6'b111111;
12'b11011110000001: data = 6'b111111;
12'b11011110000010: data = 6'b111111;
12'b11011110000011: data = 6'b111111;
12'b11011110000100: data = 6'b101010;
12'b11011110000101: data = 6'b101010;
12'b11011110000110: data = 6'b101010;
12'b11011110000111: data = 6'b101010;
12'b11011110001000: data = 6'b101010;
12'b11011110001001: data = 6'b010101;
12'b11011110001010: data = 6'b010101;
12'b11011110001011: data = 6'b010101;
12'b11011110001100: data = 6'b000000;
12'b11011110001101: data = 6'b000000;
12'b11011110001110: data = 6'b101010;
12'b11011110001111: data = 6'b101010;
12'b11011110010000: data = 6'b101010;
12'b11011110010001: data = 6'b101010;
12'b11011110010010: data = 6'b010101;
12'b11011110010011: data = 6'b010101;
12'b11011110010100: data = 6'b010101;
12'b11011110010101: data = 6'b010101;
12'b11011110010110: data = 6'b010101;
12'b11011110010111: data = 6'b010101;
12'b11011110011000: data = 6'b010101;
12'b11011110011001: data = 6'b010101;
12'b11011110011010: data = 6'b010101;
12'b11011110011011: data = 6'b010101;
12'b11011110011100: data = 6'b010101;
12'b11011110011101: data = 6'b010101;
12'b11011110011110: data = 6'b010101;
12'b11011110011111: data = 6'b010101;
12'b11011110100000: data = 6'b010101;
12'b11011110100001: data = 6'b010101;
12'b11011110100010: data = 6'b010101;
12'b11011110100011: data = 6'b010101;
12'b11011110100100: data = 6'b010101;
12'b11011110100101: data = 6'b010101;
12'b11011110100110: data = 6'b010101;
12'b11011110100111: data = 6'b010101;
12'b11011110101000: data = 6'b010101;
12'b11011110101001: data = 6'b010101;
12'b11011110101010: data = 6'b010101;
12'b111000000000: data = 6'b010101;
12'b111000000001: data = 6'b010101;
12'b111000000010: data = 6'b010101;
12'b111000000011: data = 6'b010101;
12'b111000000100: data = 6'b010101;
12'b111000000101: data = 6'b010101;
12'b111000000110: data = 6'b010101;
12'b111000000111: data = 6'b010101;
12'b111000001000: data = 6'b010101;
12'b111000001001: data = 6'b010101;
12'b111000001010: data = 6'b010101;
12'b111000001011: data = 6'b010101;
12'b111000001100: data = 6'b010101;
12'b111000001101: data = 6'b010101;
12'b111000001110: data = 6'b010101;
12'b111000001111: data = 6'b010101;
12'b111000010000: data = 6'b010101;
12'b111000010001: data = 6'b010101;
12'b111000010010: data = 6'b010101;
12'b111000010011: data = 6'b010101;
12'b111000010100: data = 6'b010101;
12'b111000010101: data = 6'b010101;
12'b111000010110: data = 6'b010101;
12'b111000010111: data = 6'b010101;
12'b111000011000: data = 6'b010101;
12'b111000011001: data = 6'b101010;
12'b111000011010: data = 6'b101010;
12'b111000011011: data = 6'b101010;
12'b111000011100: data = 6'b010101;
12'b111000011101: data = 6'b000000;
12'b111000011110: data = 6'b000000;
12'b111000011111: data = 6'b010101;
12'b111000100000: data = 6'b010101;
12'b111000100001: data = 6'b010101;
12'b111000100010: data = 6'b101010;
12'b111000100011: data = 6'b111111;
12'b111000100100: data = 6'b111111;
12'b111000100101: data = 6'b111111;
12'b111000100110: data = 6'b111111;
12'b111000100111: data = 6'b111111;
12'b111000101000: data = 6'b111111;
12'b111000101001: data = 6'b111111;
12'b111000101010: data = 6'b111111;
12'b111000101011: data = 6'b111111;
12'b111000101100: data = 6'b111111;
12'b111000101101: data = 6'b111111;
12'b111000101110: data = 6'b111111;
12'b111000101111: data = 6'b111111;
12'b111000110000: data = 6'b111111;
12'b111000110001: data = 6'b111111;
12'b111000110010: data = 6'b111111;
12'b111000110011: data = 6'b111111;
12'b111000110100: data = 6'b111111;
12'b111000110101: data = 6'b111111;
12'b111000110110: data = 6'b111111;
12'b111000110111: data = 6'b111111;
12'b111000111000: data = 6'b111111;
12'b111000111001: data = 6'b111111;
12'b111000111010: data = 6'b111111;
12'b111000111011: data = 6'b111111;
12'b111000111100: data = 6'b111111;
12'b111000111101: data = 6'b111111;
12'b111000111110: data = 6'b111111;
12'b111000111111: data = 6'b111111;
12'b1110001000000: data = 6'b111111;
12'b1110001000001: data = 6'b111111;
12'b1110001000010: data = 6'b111111;
12'b1110001000011: data = 6'b111111;
12'b1110001000100: data = 6'b111111;
12'b1110001000101: data = 6'b111111;
12'b1110001000110: data = 6'b111111;
12'b1110001000111: data = 6'b101010;
12'b1110001001000: data = 6'b101010;
12'b1110001001001: data = 6'b101010;
12'b1110001001010: data = 6'b111111;
12'b1110001001011: data = 6'b111111;
12'b1110001001100: data = 6'b111111;
12'b1110001001101: data = 6'b111111;
12'b1110001001110: data = 6'b111111;
12'b1110001001111: data = 6'b111111;
12'b1110001010000: data = 6'b111111;
12'b1110001010001: data = 6'b111111;
12'b1110001010010: data = 6'b111111;
12'b1110001010011: data = 6'b111111;
12'b1110001010100: data = 6'b111111;
12'b1110001010101: data = 6'b111111;
12'b1110001010110: data = 6'b111111;
12'b1110001010111: data = 6'b111111;
12'b1110001011000: data = 6'b111111;
12'b1110001011001: data = 6'b111111;
12'b1110001011010: data = 6'b111111;
12'b1110001011011: data = 6'b111111;
12'b1110001011100: data = 6'b111111;
12'b1110001011101: data = 6'b111111;
12'b1110001011110: data = 6'b111111;
12'b1110001011111: data = 6'b111111;
12'b1110001100000: data = 6'b111111;
12'b1110001100001: data = 6'b101010;
12'b1110001100010: data = 6'b101010;
12'b1110001100011: data = 6'b101010;
12'b1110001100100: data = 6'b111111;
12'b1110001100101: data = 6'b111111;
12'b1110001100110: data = 6'b111111;
12'b1110001100111: data = 6'b111111;
12'b1110001101000: data = 6'b111111;
12'b1110001101001: data = 6'b111111;
12'b1110001101010: data = 6'b111111;
12'b1110001101011: data = 6'b111111;
12'b1110001101100: data = 6'b111111;
12'b1110001101101: data = 6'b111111;
12'b1110001101110: data = 6'b111111;
12'b1110001101111: data = 6'b111111;
12'b1110001110000: data = 6'b111111;
12'b1110001110001: data = 6'b111111;
12'b1110001110010: data = 6'b111111;
12'b1110001110011: data = 6'b111111;
12'b1110001110100: data = 6'b111111;
12'b1110001110101: data = 6'b111111;
12'b1110001110110: data = 6'b111111;
12'b1110001110111: data = 6'b111111;
12'b1110001111000: data = 6'b111111;
12'b1110001111001: data = 6'b111111;
12'b1110001111010: data = 6'b111111;
12'b1110001111011: data = 6'b111111;
12'b1110001111100: data = 6'b111111;
12'b1110001111101: data = 6'b111111;
12'b1110001111110: data = 6'b111111;
12'b1110001111111: data = 6'b111111;
12'b11100010000000: data = 6'b111111;
12'b11100010000001: data = 6'b111111;
12'b11100010000010: data = 6'b111111;
12'b11100010000011: data = 6'b111111;
12'b11100010000100: data = 6'b111111;
12'b11100010000101: data = 6'b111111;
12'b11100010000110: data = 6'b101010;
12'b11100010000111: data = 6'b101010;
12'b11100010001000: data = 6'b101010;
12'b11100010001001: data = 6'b010101;
12'b11100010001010: data = 6'b010101;
12'b11100010001011: data = 6'b010101;
12'b11100010001100: data = 6'b000000;
12'b11100010001101: data = 6'b000000;
12'b11100010001110: data = 6'b101010;
12'b11100010001111: data = 6'b101010;
12'b11100010010000: data = 6'b101010;
12'b11100010010001: data = 6'b101010;
12'b11100010010010: data = 6'b010101;
12'b11100010010011: data = 6'b010101;
12'b11100010010100: data = 6'b010101;
12'b11100010010101: data = 6'b010101;
12'b11100010010110: data = 6'b010101;
12'b11100010010111: data = 6'b010101;
12'b11100010011000: data = 6'b010101;
12'b11100010011001: data = 6'b010101;
12'b11100010011010: data = 6'b010101;
12'b11100010011011: data = 6'b010101;
12'b11100010011100: data = 6'b010101;
12'b11100010011101: data = 6'b010101;
12'b11100010011110: data = 6'b010101;
12'b11100010011111: data = 6'b010101;
12'b11100010100000: data = 6'b010101;
12'b11100010100001: data = 6'b010101;
12'b11100010100010: data = 6'b010101;
12'b11100010100011: data = 6'b010101;
12'b11100010100100: data = 6'b010101;
12'b11100010100101: data = 6'b010101;
12'b11100010100110: data = 6'b010101;
12'b11100010100111: data = 6'b010101;
12'b11100010101000: data = 6'b010101;
12'b11100010101001: data = 6'b010101;
12'b11100010101010: data = 6'b010101;
12'b111001000000: data = 6'b010101;
12'b111001000001: data = 6'b010101;
12'b111001000010: data = 6'b010101;
12'b111001000011: data = 6'b010101;
12'b111001000100: data = 6'b010101;
12'b111001000101: data = 6'b010101;
12'b111001000110: data = 6'b010101;
12'b111001000111: data = 6'b010101;
12'b111001001000: data = 6'b010101;
12'b111001001001: data = 6'b010101;
12'b111001001010: data = 6'b010101;
12'b111001001011: data = 6'b010101;
12'b111001001100: data = 6'b010101;
12'b111001001101: data = 6'b010101;
12'b111001001110: data = 6'b010101;
12'b111001001111: data = 6'b010101;
12'b111001010000: data = 6'b010101;
12'b111001010001: data = 6'b010101;
12'b111001010010: data = 6'b010101;
12'b111001010011: data = 6'b010101;
12'b111001010100: data = 6'b010101;
12'b111001010101: data = 6'b010101;
12'b111001010110: data = 6'b010101;
12'b111001010111: data = 6'b010101;
12'b111001011000: data = 6'b010101;
12'b111001011001: data = 6'b101010;
12'b111001011010: data = 6'b101010;
12'b111001011011: data = 6'b101010;
12'b111001011100: data = 6'b010101;
12'b111001011101: data = 6'b000000;
12'b111001011110: data = 6'b000000;
12'b111001011111: data = 6'b010101;
12'b111001100000: data = 6'b010101;
12'b111001100001: data = 6'b010101;
12'b111001100010: data = 6'b101010;
12'b111001100011: data = 6'b111111;
12'b111001100100: data = 6'b111111;
12'b111001100101: data = 6'b111111;
12'b111001100110: data = 6'b111111;
12'b111001100111: data = 6'b111111;
12'b111001101000: data = 6'b111111;
12'b111001101001: data = 6'b111111;
12'b111001101010: data = 6'b111111;
12'b111001101011: data = 6'b111111;
12'b111001101100: data = 6'b111111;
12'b111001101101: data = 6'b111111;
12'b111001101110: data = 6'b111111;
12'b111001101111: data = 6'b111111;
12'b111001110000: data = 6'b111111;
12'b111001110001: data = 6'b111111;
12'b111001110010: data = 6'b111111;
12'b111001110011: data = 6'b111111;
12'b111001110100: data = 6'b111111;
12'b111001110101: data = 6'b111111;
12'b111001110110: data = 6'b111111;
12'b111001110111: data = 6'b111111;
12'b111001111000: data = 6'b111111;
12'b111001111001: data = 6'b111111;
12'b111001111010: data = 6'b111111;
12'b111001111011: data = 6'b111111;
12'b111001111100: data = 6'b111111;
12'b111001111101: data = 6'b111111;
12'b111001111110: data = 6'b111111;
12'b111001111111: data = 6'b111111;
12'b1110011000000: data = 6'b111111;
12'b1110011000001: data = 6'b111111;
12'b1110011000010: data = 6'b111111;
12'b1110011000011: data = 6'b111111;
12'b1110011000100: data = 6'b111111;
12'b1110011000101: data = 6'b111111;
12'b1110011000110: data = 6'b111111;
12'b1110011000111: data = 6'b101010;
12'b1110011001000: data = 6'b101010;
12'b1110011001001: data = 6'b101010;
12'b1110011001010: data = 6'b111111;
12'b1110011001011: data = 6'b111111;
12'b1110011001100: data = 6'b111111;
12'b1110011001101: data = 6'b111111;
12'b1110011001110: data = 6'b111111;
12'b1110011001111: data = 6'b111111;
12'b1110011010000: data = 6'b111111;
12'b1110011010001: data = 6'b111111;
12'b1110011010010: data = 6'b111111;
12'b1110011010011: data = 6'b111111;
12'b1110011010100: data = 6'b111111;
12'b1110011010101: data = 6'b111111;
12'b1110011010110: data = 6'b111111;
12'b1110011010111: data = 6'b111111;
12'b1110011011000: data = 6'b111111;
12'b1110011011001: data = 6'b111111;
12'b1110011011010: data = 6'b111111;
12'b1110011011011: data = 6'b111111;
12'b1110011011100: data = 6'b111111;
12'b1110011011101: data = 6'b111111;
12'b1110011011110: data = 6'b111111;
12'b1110011011111: data = 6'b111111;
12'b1110011100000: data = 6'b111111;
12'b1110011100001: data = 6'b101010;
12'b1110011100010: data = 6'b101010;
12'b1110011100011: data = 6'b101010;
12'b1110011100100: data = 6'b111111;
12'b1110011100101: data = 6'b111111;
12'b1110011100110: data = 6'b111111;
12'b1110011100111: data = 6'b111111;
12'b1110011101000: data = 6'b111111;
12'b1110011101001: data = 6'b111111;
12'b1110011101010: data = 6'b111111;
12'b1110011101011: data = 6'b111111;
12'b1110011101100: data = 6'b111111;
12'b1110011101101: data = 6'b111111;
12'b1110011101110: data = 6'b111111;
12'b1110011101111: data = 6'b111111;
12'b1110011110000: data = 6'b111111;
12'b1110011110001: data = 6'b111111;
12'b1110011110010: data = 6'b111111;
12'b1110011110011: data = 6'b111111;
12'b1110011110100: data = 6'b111111;
12'b1110011110101: data = 6'b111111;
12'b1110011110110: data = 6'b111111;
12'b1110011110111: data = 6'b111111;
12'b1110011111000: data = 6'b111111;
12'b1110011111001: data = 6'b111111;
12'b1110011111010: data = 6'b111111;
12'b1110011111011: data = 6'b111111;
12'b1110011111100: data = 6'b111111;
12'b1110011111101: data = 6'b111111;
12'b1110011111110: data = 6'b111111;
12'b1110011111111: data = 6'b111111;
12'b11100110000000: data = 6'b111111;
12'b11100110000001: data = 6'b111111;
12'b11100110000010: data = 6'b111111;
12'b11100110000011: data = 6'b111111;
12'b11100110000100: data = 6'b111111;
12'b11100110000101: data = 6'b111111;
12'b11100110000110: data = 6'b111111;
12'b11100110000111: data = 6'b111111;
12'b11100110001000: data = 6'b101010;
12'b11100110001001: data = 6'b010101;
12'b11100110001010: data = 6'b010101;
12'b11100110001011: data = 6'b010101;
12'b11100110001100: data = 6'b000000;
12'b11100110001101: data = 6'b000000;
12'b11100110001110: data = 6'b101010;
12'b11100110001111: data = 6'b101010;
12'b11100110010000: data = 6'b101010;
12'b11100110010001: data = 6'b101010;
12'b11100110010010: data = 6'b010101;
12'b11100110010011: data = 6'b010101;
12'b11100110010100: data = 6'b010101;
12'b11100110010101: data = 6'b010101;
12'b11100110010110: data = 6'b010101;
12'b11100110010111: data = 6'b010101;
12'b11100110011000: data = 6'b010101;
12'b11100110011001: data = 6'b010101;
12'b11100110011010: data = 6'b010101;
12'b11100110011011: data = 6'b010101;
12'b11100110011100: data = 6'b010101;
12'b11100110011101: data = 6'b010101;
12'b11100110011110: data = 6'b010101;
12'b11100110011111: data = 6'b010101;
12'b11100110100000: data = 6'b010101;
12'b11100110100001: data = 6'b010101;
12'b11100110100010: data = 6'b010101;
12'b11100110100011: data = 6'b010101;
12'b11100110100100: data = 6'b010101;
12'b11100110100101: data = 6'b010101;
12'b11100110100110: data = 6'b010101;
12'b11100110100111: data = 6'b010101;
12'b11100110101000: data = 6'b010101;
12'b11100110101001: data = 6'b010101;
12'b11100110101010: data = 6'b010101;
12'b111010000000: data = 6'b010101;
12'b111010000001: data = 6'b010101;
12'b111010000010: data = 6'b010101;
12'b111010000011: data = 6'b010101;
12'b111010000100: data = 6'b010101;
12'b111010000101: data = 6'b010101;
12'b111010000110: data = 6'b010101;
12'b111010000111: data = 6'b010101;
12'b111010001000: data = 6'b010101;
12'b111010001001: data = 6'b010101;
12'b111010001010: data = 6'b010101;
12'b111010001011: data = 6'b010101;
12'b111010001100: data = 6'b010101;
12'b111010001101: data = 6'b010101;
12'b111010001110: data = 6'b010101;
12'b111010001111: data = 6'b010101;
12'b111010010000: data = 6'b010101;
12'b111010010001: data = 6'b010101;
12'b111010010010: data = 6'b010101;
12'b111010010011: data = 6'b010101;
12'b111010010100: data = 6'b010101;
12'b111010010101: data = 6'b010101;
12'b111010010110: data = 6'b010101;
12'b111010010111: data = 6'b010101;
12'b111010011000: data = 6'b010101;
12'b111010011001: data = 6'b101010;
12'b111010011010: data = 6'b101010;
12'b111010011011: data = 6'b101010;
12'b111010011100: data = 6'b010101;
12'b111010011101: data = 6'b000000;
12'b111010011110: data = 6'b000000;
12'b111010011111: data = 6'b010101;
12'b111010100000: data = 6'b010101;
12'b111010100001: data = 6'b010101;
12'b111010100010: data = 6'b101010;
12'b111010100011: data = 6'b111111;
12'b111010100100: data = 6'b111111;
12'b111010100101: data = 6'b111111;
12'b111010100110: data = 6'b111111;
12'b111010100111: data = 6'b111111;
12'b111010101000: data = 6'b111111;
12'b111010101001: data = 6'b111111;
12'b111010101010: data = 6'b111111;
12'b111010101011: data = 6'b111111;
12'b111010101100: data = 6'b111111;
12'b111010101101: data = 6'b111111;
12'b111010101110: data = 6'b111111;
12'b111010101111: data = 6'b111111;
12'b111010110000: data = 6'b111111;
12'b111010110001: data = 6'b111111;
12'b111010110010: data = 6'b111111;
12'b111010110011: data = 6'b111111;
12'b111010110100: data = 6'b111111;
12'b111010110101: data = 6'b111111;
12'b111010110110: data = 6'b111111;
12'b111010110111: data = 6'b111111;
12'b111010111000: data = 6'b111111;
12'b111010111001: data = 6'b111111;
12'b111010111010: data = 6'b111111;
12'b111010111011: data = 6'b111111;
12'b111010111100: data = 6'b111111;
12'b111010111101: data = 6'b111111;
12'b111010111110: data = 6'b111111;
12'b111010111111: data = 6'b111111;
12'b1110101000000: data = 6'b111111;
12'b1110101000001: data = 6'b111111;
12'b1110101000010: data = 6'b111111;
12'b1110101000011: data = 6'b111111;
12'b1110101000100: data = 6'b111111;
12'b1110101000101: data = 6'b111111;
12'b1110101000110: data = 6'b111111;
12'b1110101000111: data = 6'b101010;
12'b1110101001000: data = 6'b101010;
12'b1110101001001: data = 6'b101010;
12'b1110101001010: data = 6'b111111;
12'b1110101001011: data = 6'b111111;
12'b1110101001100: data = 6'b111111;
12'b1110101001101: data = 6'b111111;
12'b1110101001110: data = 6'b111111;
12'b1110101001111: data = 6'b111111;
12'b1110101010000: data = 6'b111111;
12'b1110101010001: data = 6'b111111;
12'b1110101010010: data = 6'b111111;
12'b1110101010011: data = 6'b111111;
12'b1110101010100: data = 6'b111111;
12'b1110101010101: data = 6'b111111;
12'b1110101010110: data = 6'b111111;
12'b1110101010111: data = 6'b111111;
12'b1110101011000: data = 6'b111111;
12'b1110101011001: data = 6'b111111;
12'b1110101011010: data = 6'b111111;
12'b1110101011011: data = 6'b111111;
12'b1110101011100: data = 6'b111111;
12'b1110101011101: data = 6'b111111;
12'b1110101011110: data = 6'b111111;
12'b1110101011111: data = 6'b111111;
12'b1110101100000: data = 6'b111111;
12'b1110101100001: data = 6'b101010;
12'b1110101100010: data = 6'b101010;
12'b1110101100011: data = 6'b101010;
12'b1110101100100: data = 6'b111111;
12'b1110101100101: data = 6'b111111;
12'b1110101100110: data = 6'b111111;
12'b1110101100111: data = 6'b111111;
12'b1110101101000: data = 6'b111111;
12'b1110101101001: data = 6'b111111;
12'b1110101101010: data = 6'b111111;
12'b1110101101011: data = 6'b111111;
12'b1110101101100: data = 6'b111111;
12'b1110101101101: data = 6'b111111;
12'b1110101101110: data = 6'b111111;
12'b1110101101111: data = 6'b111111;
12'b1110101110000: data = 6'b111111;
12'b1110101110001: data = 6'b111111;
12'b1110101110010: data = 6'b111111;
12'b1110101110011: data = 6'b111111;
12'b1110101110100: data = 6'b111111;
12'b1110101110101: data = 6'b111111;
12'b1110101110110: data = 6'b111111;
12'b1110101110111: data = 6'b111111;
12'b1110101111000: data = 6'b111111;
12'b1110101111001: data = 6'b111111;
12'b1110101111010: data = 6'b111111;
12'b1110101111011: data = 6'b111111;
12'b1110101111100: data = 6'b111111;
12'b1110101111101: data = 6'b111111;
12'b1110101111110: data = 6'b111111;
12'b1110101111111: data = 6'b111111;
12'b11101010000000: data = 6'b111111;
12'b11101010000001: data = 6'b111111;
12'b11101010000010: data = 6'b111111;
12'b11101010000011: data = 6'b111111;
12'b11101010000100: data = 6'b111111;
12'b11101010000101: data = 6'b111111;
12'b11101010000110: data = 6'b111111;
12'b11101010000111: data = 6'b111111;
12'b11101010001000: data = 6'b101010;
12'b11101010001001: data = 6'b010101;
12'b11101010001010: data = 6'b010101;
12'b11101010001011: data = 6'b010101;
12'b11101010001100: data = 6'b000000;
12'b11101010001101: data = 6'b000000;
12'b11101010001110: data = 6'b101010;
12'b11101010001111: data = 6'b101010;
12'b11101010010000: data = 6'b101010;
12'b11101010010001: data = 6'b101010;
12'b11101010010010: data = 6'b010101;
12'b11101010010011: data = 6'b010101;
12'b11101010010100: data = 6'b010101;
12'b11101010010101: data = 6'b010101;
12'b11101010010110: data = 6'b010101;
12'b11101010010111: data = 6'b010101;
12'b11101010011000: data = 6'b010101;
12'b11101010011001: data = 6'b010101;
12'b11101010011010: data = 6'b010101;
12'b11101010011011: data = 6'b010101;
12'b11101010011100: data = 6'b010101;
12'b11101010011101: data = 6'b010101;
12'b11101010011110: data = 6'b010101;
12'b11101010011111: data = 6'b010101;
12'b11101010100000: data = 6'b010101;
12'b11101010100001: data = 6'b010101;
12'b11101010100010: data = 6'b010101;
12'b11101010100011: data = 6'b010101;
12'b11101010100100: data = 6'b010101;
12'b11101010100101: data = 6'b010101;
12'b11101010100110: data = 6'b010101;
12'b11101010100111: data = 6'b010101;
12'b11101010101000: data = 6'b010101;
12'b11101010101001: data = 6'b010101;
12'b11101010101010: data = 6'b010101;
12'b111011000000: data = 6'b010101;
12'b111011000001: data = 6'b010101;
12'b111011000010: data = 6'b010101;
12'b111011000011: data = 6'b010101;
12'b111011000100: data = 6'b010101;
12'b111011000101: data = 6'b010101;
12'b111011000110: data = 6'b010101;
12'b111011000111: data = 6'b010101;
12'b111011001000: data = 6'b010101;
12'b111011001001: data = 6'b010101;
12'b111011001010: data = 6'b010101;
12'b111011001011: data = 6'b010101;
12'b111011001100: data = 6'b010101;
12'b111011001101: data = 6'b010101;
12'b111011001110: data = 6'b010101;
12'b111011001111: data = 6'b010101;
12'b111011010000: data = 6'b010101;
12'b111011010001: data = 6'b010101;
12'b111011010010: data = 6'b010101;
12'b111011010011: data = 6'b010101;
12'b111011010100: data = 6'b010101;
12'b111011010101: data = 6'b010101;
12'b111011010110: data = 6'b010101;
12'b111011010111: data = 6'b010101;
12'b111011011000: data = 6'b010101;
12'b111011011001: data = 6'b101010;
12'b111011011010: data = 6'b101010;
12'b111011011011: data = 6'b101010;
12'b111011011100: data = 6'b010101;
12'b111011011101: data = 6'b000000;
12'b111011011110: data = 6'b000000;
12'b111011011111: data = 6'b010101;
12'b111011100000: data = 6'b010101;
12'b111011100001: data = 6'b010101;
12'b111011100010: data = 6'b101010;
12'b111011100011: data = 6'b111111;
12'b111011100100: data = 6'b111111;
12'b111011100101: data = 6'b111111;
12'b111011100110: data = 6'b111111;
12'b111011100111: data = 6'b111111;
12'b111011101000: data = 6'b111111;
12'b111011101001: data = 6'b111111;
12'b111011101010: data = 6'b111111;
12'b111011101011: data = 6'b111111;
12'b111011101100: data = 6'b111111;
12'b111011101101: data = 6'b111111;
12'b111011101110: data = 6'b111111;
12'b111011101111: data = 6'b111111;
12'b111011110000: data = 6'b111111;
12'b111011110001: data = 6'b111111;
12'b111011110010: data = 6'b111111;
12'b111011110011: data = 6'b111111;
12'b111011110100: data = 6'b111111;
12'b111011110101: data = 6'b111111;
12'b111011110110: data = 6'b111111;
12'b111011110111: data = 6'b111111;
12'b111011111000: data = 6'b111111;
12'b111011111001: data = 6'b111111;
12'b111011111010: data = 6'b111111;
12'b111011111011: data = 6'b111111;
12'b111011111100: data = 6'b111111;
12'b111011111101: data = 6'b111111;
12'b111011111110: data = 6'b111111;
12'b111011111111: data = 6'b111111;
12'b1110111000000: data = 6'b111111;
12'b1110111000001: data = 6'b111111;
12'b1110111000010: data = 6'b111111;
12'b1110111000011: data = 6'b111111;
12'b1110111000100: data = 6'b111111;
12'b1110111000101: data = 6'b111111;
12'b1110111000110: data = 6'b111111;
12'b1110111000111: data = 6'b101010;
12'b1110111001000: data = 6'b101010;
12'b1110111001001: data = 6'b101010;
12'b1110111001010: data = 6'b111111;
12'b1110111001011: data = 6'b111111;
12'b1110111001100: data = 6'b111111;
12'b1110111001101: data = 6'b111111;
12'b1110111001110: data = 6'b111111;
12'b1110111001111: data = 6'b111111;
12'b1110111010000: data = 6'b111111;
12'b1110111010001: data = 6'b111111;
12'b1110111010010: data = 6'b111111;
12'b1110111010011: data = 6'b111111;
12'b1110111010100: data = 6'b111111;
12'b1110111010101: data = 6'b111111;
12'b1110111010110: data = 6'b111111;
12'b1110111010111: data = 6'b111111;
12'b1110111011000: data = 6'b111111;
12'b1110111011001: data = 6'b111111;
12'b1110111011010: data = 6'b111111;
12'b1110111011011: data = 6'b111111;
12'b1110111011100: data = 6'b111111;
12'b1110111011101: data = 6'b111111;
12'b1110111011110: data = 6'b111111;
12'b1110111011111: data = 6'b111111;
12'b1110111100000: data = 6'b111111;
12'b1110111100001: data = 6'b101010;
12'b1110111100010: data = 6'b101010;
12'b1110111100011: data = 6'b101010;
12'b1110111100100: data = 6'b111111;
12'b1110111100101: data = 6'b111111;
12'b1110111100110: data = 6'b111111;
12'b1110111100111: data = 6'b111111;
12'b1110111101000: data = 6'b111111;
12'b1110111101001: data = 6'b111111;
12'b1110111101010: data = 6'b111111;
12'b1110111101011: data = 6'b111111;
12'b1110111101100: data = 6'b111111;
12'b1110111101101: data = 6'b111111;
12'b1110111101110: data = 6'b111111;
12'b1110111101111: data = 6'b111111;
12'b1110111110000: data = 6'b111111;
12'b1110111110001: data = 6'b111111;
12'b1110111110010: data = 6'b111111;
12'b1110111110011: data = 6'b111111;
12'b1110111110100: data = 6'b111111;
12'b1110111110101: data = 6'b111111;
12'b1110111110110: data = 6'b111111;
12'b1110111110111: data = 6'b111111;
12'b1110111111000: data = 6'b111111;
12'b1110111111001: data = 6'b111111;
12'b1110111111010: data = 6'b111111;
12'b1110111111011: data = 6'b111111;
12'b1110111111100: data = 6'b111111;
12'b1110111111101: data = 6'b111111;
12'b1110111111110: data = 6'b111111;
12'b1110111111111: data = 6'b111111;
12'b11101110000000: data = 6'b111111;
12'b11101110000001: data = 6'b111111;
12'b11101110000010: data = 6'b111111;
12'b11101110000011: data = 6'b111111;
12'b11101110000100: data = 6'b111111;
12'b11101110000101: data = 6'b111111;
12'b11101110000110: data = 6'b111111;
12'b11101110000111: data = 6'b111111;
12'b11101110001000: data = 6'b101010;
12'b11101110001001: data = 6'b010101;
12'b11101110001010: data = 6'b010101;
12'b11101110001011: data = 6'b010101;
12'b11101110001100: data = 6'b000000;
12'b11101110001101: data = 6'b000000;
12'b11101110001110: data = 6'b101010;
12'b11101110001111: data = 6'b101010;
12'b11101110010000: data = 6'b101010;
12'b11101110010001: data = 6'b101010;
12'b11101110010010: data = 6'b010101;
12'b11101110010011: data = 6'b010101;
12'b11101110010100: data = 6'b010101;
12'b11101110010101: data = 6'b010101;
12'b11101110010110: data = 6'b010101;
12'b11101110010111: data = 6'b010101;
12'b11101110011000: data = 6'b010101;
12'b11101110011001: data = 6'b010101;
12'b11101110011010: data = 6'b010101;
12'b11101110011011: data = 6'b010101;
12'b11101110011100: data = 6'b010101;
12'b11101110011101: data = 6'b010101;
12'b11101110011110: data = 6'b010101;
12'b11101110011111: data = 6'b010101;
12'b11101110100000: data = 6'b010101;
12'b11101110100001: data = 6'b010101;
12'b11101110100010: data = 6'b010101;
12'b11101110100011: data = 6'b010101;
12'b11101110100100: data = 6'b010101;
12'b11101110100101: data = 6'b010101;
12'b11101110100110: data = 6'b010101;
12'b11101110100111: data = 6'b010101;
12'b11101110101000: data = 6'b010101;
12'b11101110101001: data = 6'b010101;
12'b11101110101010: data = 6'b010101;
12'b111100000000: data = 6'b010101;
12'b111100000001: data = 6'b010101;
12'b111100000010: data = 6'b010101;
12'b111100000011: data = 6'b010101;
12'b111100000100: data = 6'b010101;
12'b111100000101: data = 6'b010101;
12'b111100000110: data = 6'b010101;
12'b111100000111: data = 6'b010101;
12'b111100001000: data = 6'b010101;
12'b111100001001: data = 6'b010101;
12'b111100001010: data = 6'b010101;
12'b111100001011: data = 6'b010101;
12'b111100001100: data = 6'b010101;
12'b111100001101: data = 6'b010101;
12'b111100001110: data = 6'b010101;
12'b111100001111: data = 6'b010101;
12'b111100010000: data = 6'b010101;
12'b111100010001: data = 6'b010101;
12'b111100010010: data = 6'b010101;
12'b111100010011: data = 6'b010101;
12'b111100010100: data = 6'b010101;
12'b111100010101: data = 6'b010101;
12'b111100010110: data = 6'b010101;
12'b111100010111: data = 6'b010101;
12'b111100011000: data = 6'b010101;
12'b111100011001: data = 6'b101010;
12'b111100011010: data = 6'b101010;
12'b111100011011: data = 6'b101010;
12'b111100011100: data = 6'b010101;
12'b111100011101: data = 6'b000000;
12'b111100011110: data = 6'b000000;
12'b111100011111: data = 6'b010101;
12'b111100100000: data = 6'b010101;
12'b111100100001: data = 6'b010101;
12'b111100100010: data = 6'b101010;
12'b111100100011: data = 6'b111111;
12'b111100100100: data = 6'b111111;
12'b111100100101: data = 6'b111111;
12'b111100100110: data = 6'b111111;
12'b111100100111: data = 6'b111111;
12'b111100101000: data = 6'b111111;
12'b111100101001: data = 6'b111111;
12'b111100101010: data = 6'b111111;
12'b111100101011: data = 6'b111111;
12'b111100101100: data = 6'b111111;
12'b111100101101: data = 6'b111111;
12'b111100101110: data = 6'b111111;
12'b111100101111: data = 6'b111111;
12'b111100110000: data = 6'b111111;
12'b111100110001: data = 6'b111111;
12'b111100110010: data = 6'b111111;
12'b111100110011: data = 6'b111111;
12'b111100110100: data = 6'b111111;
12'b111100110101: data = 6'b111111;
12'b111100110110: data = 6'b111111;
12'b111100110111: data = 6'b111111;
12'b111100111000: data = 6'b111111;
12'b111100111001: data = 6'b111111;
12'b111100111010: data = 6'b111111;
12'b111100111011: data = 6'b111111;
12'b111100111100: data = 6'b111111;
12'b111100111101: data = 6'b111111;
12'b111100111110: data = 6'b111111;
12'b111100111111: data = 6'b111111;
12'b1111001000000: data = 6'b111111;
12'b1111001000001: data = 6'b111111;
12'b1111001000010: data = 6'b111111;
12'b1111001000011: data = 6'b111111;
12'b1111001000100: data = 6'b111111;
12'b1111001000101: data = 6'b111111;
12'b1111001000110: data = 6'b111111;
12'b1111001000111: data = 6'b101010;
12'b1111001001000: data = 6'b101010;
12'b1111001001001: data = 6'b101010;
12'b1111001001010: data = 6'b111111;
12'b1111001001011: data = 6'b111111;
12'b1111001001100: data = 6'b111111;
12'b1111001001101: data = 6'b111111;
12'b1111001001110: data = 6'b111111;
12'b1111001001111: data = 6'b111111;
12'b1111001010000: data = 6'b111111;
12'b1111001010001: data = 6'b111111;
12'b1111001010010: data = 6'b111111;
12'b1111001010011: data = 6'b111111;
12'b1111001010100: data = 6'b111111;
12'b1111001010101: data = 6'b111111;
12'b1111001010110: data = 6'b111111;
12'b1111001010111: data = 6'b111111;
12'b1111001011000: data = 6'b111111;
12'b1111001011001: data = 6'b111111;
12'b1111001011010: data = 6'b111111;
12'b1111001011011: data = 6'b111111;
12'b1111001011100: data = 6'b111111;
12'b1111001011101: data = 6'b111111;
12'b1111001011110: data = 6'b111111;
12'b1111001011111: data = 6'b111111;
12'b1111001100000: data = 6'b111111;
12'b1111001100001: data = 6'b101010;
12'b1111001100010: data = 6'b101010;
12'b1111001100011: data = 6'b101010;
12'b1111001100100: data = 6'b111111;
12'b1111001100101: data = 6'b111111;
12'b1111001100110: data = 6'b111111;
12'b1111001100111: data = 6'b111111;
12'b1111001101000: data = 6'b111111;
12'b1111001101001: data = 6'b111111;
12'b1111001101010: data = 6'b111111;
12'b1111001101011: data = 6'b111111;
12'b1111001101100: data = 6'b111111;
12'b1111001101101: data = 6'b111111;
12'b1111001101110: data = 6'b111111;
12'b1111001101111: data = 6'b111111;
12'b1111001110000: data = 6'b111111;
12'b1111001110001: data = 6'b111111;
12'b1111001110010: data = 6'b111111;
12'b1111001110011: data = 6'b111111;
12'b1111001110100: data = 6'b111111;
12'b1111001110101: data = 6'b111111;
12'b1111001110110: data = 6'b111111;
12'b1111001110111: data = 6'b111111;
12'b1111001111000: data = 6'b111111;
12'b1111001111001: data = 6'b111111;
12'b1111001111010: data = 6'b111111;
12'b1111001111011: data = 6'b111111;
12'b1111001111100: data = 6'b111111;
12'b1111001111101: data = 6'b111111;
12'b1111001111110: data = 6'b111111;
12'b1111001111111: data = 6'b111111;
12'b11110010000000: data = 6'b111111;
12'b11110010000001: data = 6'b111111;
12'b11110010000010: data = 6'b111111;
12'b11110010000011: data = 6'b111111;
12'b11110010000100: data = 6'b111111;
12'b11110010000101: data = 6'b111111;
12'b11110010000110: data = 6'b111111;
12'b11110010000111: data = 6'b111111;
12'b11110010001000: data = 6'b101010;
12'b11110010001001: data = 6'b010101;
12'b11110010001010: data = 6'b010101;
12'b11110010001011: data = 6'b010101;
12'b11110010001100: data = 6'b000000;
12'b11110010001101: data = 6'b000000;
12'b11110010001110: data = 6'b101010;
12'b11110010001111: data = 6'b101010;
12'b11110010010000: data = 6'b101010;
12'b11110010010001: data = 6'b101010;
12'b11110010010010: data = 6'b010101;
12'b11110010010011: data = 6'b010101;
12'b11110010010100: data = 6'b010101;
12'b11110010010101: data = 6'b010101;
12'b11110010010110: data = 6'b010101;
12'b11110010010111: data = 6'b010101;
12'b11110010011000: data = 6'b010101;
12'b11110010011001: data = 6'b010101;
12'b11110010011010: data = 6'b010101;
12'b11110010011011: data = 6'b010101;
12'b11110010011100: data = 6'b010101;
12'b11110010011101: data = 6'b010101;
12'b11110010011110: data = 6'b010101;
12'b11110010011111: data = 6'b010101;
12'b11110010100000: data = 6'b010101;
12'b11110010100001: data = 6'b010101;
12'b11110010100010: data = 6'b010101;
12'b11110010100011: data = 6'b010101;
12'b11110010100100: data = 6'b010101;
12'b11110010100101: data = 6'b010101;
12'b11110010100110: data = 6'b010101;
12'b11110010100111: data = 6'b010101;
12'b11110010101000: data = 6'b010101;
12'b11110010101001: data = 6'b010101;
12'b11110010101010: data = 6'b010101;
12'b111101000000: data = 6'b010101;
12'b111101000001: data = 6'b010101;
12'b111101000010: data = 6'b010101;
12'b111101000011: data = 6'b010101;
12'b111101000100: data = 6'b010101;
12'b111101000101: data = 6'b010101;
12'b111101000110: data = 6'b010101;
12'b111101000111: data = 6'b010101;
12'b111101001000: data = 6'b010101;
12'b111101001001: data = 6'b010101;
12'b111101001010: data = 6'b010101;
12'b111101001011: data = 6'b010101;
12'b111101001100: data = 6'b010101;
12'b111101001101: data = 6'b010101;
12'b111101001110: data = 6'b010101;
12'b111101001111: data = 6'b010101;
12'b111101010000: data = 6'b010101;
12'b111101010001: data = 6'b010101;
12'b111101010010: data = 6'b010101;
12'b111101010011: data = 6'b010101;
12'b111101010100: data = 6'b010101;
12'b111101010101: data = 6'b010101;
12'b111101010110: data = 6'b010101;
12'b111101010111: data = 6'b010101;
12'b111101011000: data = 6'b010101;
12'b111101011001: data = 6'b101010;
12'b111101011010: data = 6'b101010;
12'b111101011011: data = 6'b101010;
12'b111101011100: data = 6'b010101;
12'b111101011101: data = 6'b000000;
12'b111101011110: data = 6'b000000;
12'b111101011111: data = 6'b010101;
12'b111101100000: data = 6'b010101;
12'b111101100001: data = 6'b010101;
12'b111101100010: data = 6'b101010;
12'b111101100011: data = 6'b101010;
12'b111101100100: data = 6'b101010;
12'b111101100101: data = 6'b111110;
12'b111101100110: data = 6'b111110;
12'b111101100111: data = 6'b111111;
12'b111101101000: data = 6'b111111;
12'b111101101001: data = 6'b111111;
12'b111101101010: data = 6'b111111;
12'b111101101011: data = 6'b111111;
12'b111101101100: data = 6'b111111;
12'b111101101101: data = 6'b111111;
12'b111101101110: data = 6'b111111;
12'b111101101111: data = 6'b111111;
12'b111101110000: data = 6'b111111;
12'b111101110001: data = 6'b111111;
12'b111101110010: data = 6'b111111;
12'b111101110011: data = 6'b111111;
12'b111101110100: data = 6'b111111;
12'b111101110101: data = 6'b111111;
12'b111101110110: data = 6'b111111;
12'b111101110111: data = 6'b111111;
12'b111101111000: data = 6'b111111;
12'b111101111001: data = 6'b111111;
12'b111101111010: data = 6'b111111;
12'b111101111011: data = 6'b111111;
12'b111101111100: data = 6'b111111;
12'b111101111101: data = 6'b111111;
12'b111101111110: data = 6'b111111;
12'b111101111111: data = 6'b111111;
12'b1111011000000: data = 6'b111111;
12'b1111011000001: data = 6'b111111;
12'b1111011000010: data = 6'b101010;
12'b1111011000011: data = 6'b101010;
12'b1111011000100: data = 6'b111110;
12'b1111011000101: data = 6'b111111;
12'b1111011000110: data = 6'b111111;
12'b1111011000111: data = 6'b101010;
12'b1111011001000: data = 6'b101010;
12'b1111011001001: data = 6'b101010;
12'b1111011001010: data = 6'b111111;
12'b1111011001011: data = 6'b111111;
12'b1111011001100: data = 6'b111111;
12'b1111011001101: data = 6'b111111;
12'b1111011001110: data = 6'b111111;
12'b1111011001111: data = 6'b111111;
12'b1111011010000: data = 6'b111111;
12'b1111011010001: data = 6'b111111;
12'b1111011010010: data = 6'b111111;
12'b1111011010011: data = 6'b111111;
12'b1111011010100: data = 6'b111111;
12'b1111011010101: data = 6'b111111;
12'b1111011010110: data = 6'b111111;
12'b1111011010111: data = 6'b111111;
12'b1111011011000: data = 6'b111111;
12'b1111011011001: data = 6'b111111;
12'b1111011011010: data = 6'b111111;
12'b1111011011011: data = 6'b111111;
12'b1111011011100: data = 6'b111111;
12'b1111011011101: data = 6'b111111;
12'b1111011011110: data = 6'b111111;
12'b1111011011111: data = 6'b111111;
12'b1111011100000: data = 6'b111111;
12'b1111011100001: data = 6'b101010;
12'b1111011100010: data = 6'b101010;
12'b1111011100011: data = 6'b101010;
12'b1111011100100: data = 6'b111111;
12'b1111011100101: data = 6'b111111;
12'b1111011100110: data = 6'b111111;
12'b1111011100111: data = 6'b111111;
12'b1111011101000: data = 6'b111111;
12'b1111011101001: data = 6'b111111;
12'b1111011101010: data = 6'b111111;
12'b1111011101011: data = 6'b111111;
12'b1111011101100: data = 6'b111111;
12'b1111011101101: data = 6'b111111;
12'b1111011101110: data = 6'b111111;
12'b1111011101111: data = 6'b111111;
12'b1111011110000: data = 6'b111111;
12'b1111011110001: data = 6'b111111;
12'b1111011110010: data = 6'b111111;
12'b1111011110011: data = 6'b111111;
12'b1111011110100: data = 6'b111111;
12'b1111011110101: data = 6'b111111;
12'b1111011110110: data = 6'b111111;
12'b1111011110111: data = 6'b111111;
12'b1111011111000: data = 6'b111111;
12'b1111011111001: data = 6'b111111;
12'b1111011111010: data = 6'b111111;
12'b1111011111011: data = 6'b111111;
12'b1111011111100: data = 6'b111111;
12'b1111011111101: data = 6'b111111;
12'b1111011111110: data = 6'b111111;
12'b1111011111111: data = 6'b111111;
12'b11110110000000: data = 6'b111111;
12'b11110110000001: data = 6'b111111;
12'b11110110000010: data = 6'b111111;
12'b11110110000011: data = 6'b111111;
12'b11110110000100: data = 6'b111111;
12'b11110110000101: data = 6'b111111;
12'b11110110000110: data = 6'b111110;
12'b11110110000111: data = 6'b111110;
12'b11110110001000: data = 6'b101010;
12'b11110110001001: data = 6'b010101;
12'b11110110001010: data = 6'b010101;
12'b11110110001011: data = 6'b010101;
12'b11110110001100: data = 6'b000000;
12'b11110110001101: data = 6'b000000;
12'b11110110001110: data = 6'b101010;
12'b11110110001111: data = 6'b101010;
12'b11110110010000: data = 6'b101010;
12'b11110110010001: data = 6'b101010;
12'b11110110010010: data = 6'b010101;
12'b11110110010011: data = 6'b010101;
12'b11110110010100: data = 6'b010101;
12'b11110110010101: data = 6'b010101;
12'b11110110010110: data = 6'b010101;
12'b11110110010111: data = 6'b010101;
12'b11110110011000: data = 6'b010101;
12'b11110110011001: data = 6'b010101;
12'b11110110011010: data = 6'b010101;
12'b11110110011011: data = 6'b010101;
12'b11110110011100: data = 6'b010101;
12'b11110110011101: data = 6'b010101;
12'b11110110011110: data = 6'b010101;
12'b11110110011111: data = 6'b010101;
12'b11110110100000: data = 6'b010101;
12'b11110110100001: data = 6'b010101;
12'b11110110100010: data = 6'b010101;
12'b11110110100011: data = 6'b010101;
12'b11110110100100: data = 6'b010101;
12'b11110110100101: data = 6'b010101;
12'b11110110100110: data = 6'b010101;
12'b11110110100111: data = 6'b010101;
12'b11110110101000: data = 6'b010101;
12'b11110110101001: data = 6'b010101;
12'b11110110101010: data = 6'b010101;
12'b111110000000: data = 6'b010101;
12'b111110000001: data = 6'b010101;
12'b111110000010: data = 6'b010101;
12'b111110000011: data = 6'b010101;
12'b111110000100: data = 6'b010101;
12'b111110000101: data = 6'b010101;
12'b111110000110: data = 6'b010101;
12'b111110000111: data = 6'b010101;
12'b111110001000: data = 6'b010101;
12'b111110001001: data = 6'b010101;
12'b111110001010: data = 6'b010101;
12'b111110001011: data = 6'b010101;
12'b111110001100: data = 6'b010101;
12'b111110001101: data = 6'b010101;
12'b111110001110: data = 6'b010101;
12'b111110001111: data = 6'b010101;
12'b111110010000: data = 6'b010101;
12'b111110010001: data = 6'b010101;
12'b111110010010: data = 6'b010101;
12'b111110010011: data = 6'b010101;
12'b111110010100: data = 6'b010101;
12'b111110010101: data = 6'b010101;
12'b111110010110: data = 6'b010101;
12'b111110010111: data = 6'b010101;
12'b111110011000: data = 6'b010101;
12'b111110011001: data = 6'b101010;
12'b111110011010: data = 6'b101010;
12'b111110011011: data = 6'b101010;
12'b111110011100: data = 6'b010101;
12'b111110011101: data = 6'b000000;
12'b111110011110: data = 6'b000000;
12'b111110011111: data = 6'b010101;
12'b111110100000: data = 6'b010101;
12'b111110100001: data = 6'b010101;
12'b111110100010: data = 6'b101010;
12'b111110100011: data = 6'b101010;
12'b111110100100: data = 6'b101010;
12'b111110100101: data = 6'b111010;
12'b111110100110: data = 6'b111110;
12'b111110100111: data = 6'b111111;
12'b111110101000: data = 6'b111111;
12'b111110101001: data = 6'b111111;
12'b111110101010: data = 6'b111111;
12'b111110101011: data = 6'b111111;
12'b111110101100: data = 6'b111111;
12'b111110101101: data = 6'b111111;
12'b111110101110: data = 6'b111111;
12'b111110101111: data = 6'b111111;
12'b111110110000: data = 6'b111111;
12'b111110110001: data = 6'b111111;
12'b111110110010: data = 6'b111111;
12'b111110110011: data = 6'b111111;
12'b111110110100: data = 6'b111111;
12'b111110110101: data = 6'b111111;
12'b111110110110: data = 6'b111111;
12'b111110110111: data = 6'b111111;
12'b111110111000: data = 6'b111111;
12'b111110111001: data = 6'b111111;
12'b111110111010: data = 6'b111111;
12'b111110111011: data = 6'b111111;
12'b111110111100: data = 6'b111111;
12'b111110111101: data = 6'b111111;
12'b111110111110: data = 6'b111111;
12'b111110111111: data = 6'b111111;
12'b1111101000000: data = 6'b111111;
12'b1111101000001: data = 6'b111110;
12'b1111101000010: data = 6'b101010;
12'b1111101000011: data = 6'b101010;
12'b1111101000100: data = 6'b101010;
12'b1111101000101: data = 6'b111111;
12'b1111101000110: data = 6'b111111;
12'b1111101000111: data = 6'b101010;
12'b1111101001000: data = 6'b101010;
12'b1111101001001: data = 6'b101010;
12'b1111101001010: data = 6'b111111;
12'b1111101001011: data = 6'b111111;
12'b1111101001100: data = 6'b111111;
12'b1111101001101: data = 6'b111111;
12'b1111101001110: data = 6'b111111;
12'b1111101001111: data = 6'b111111;
12'b1111101010000: data = 6'b111111;
12'b1111101010001: data = 6'b111111;
12'b1111101010010: data = 6'b111111;
12'b1111101010011: data = 6'b111111;
12'b1111101010100: data = 6'b111111;
12'b1111101010101: data = 6'b111111;
12'b1111101010110: data = 6'b111111;
12'b1111101010111: data = 6'b111111;
12'b1111101011000: data = 6'b111111;
12'b1111101011001: data = 6'b111111;
12'b1111101011010: data = 6'b111111;
12'b1111101011011: data = 6'b111111;
12'b1111101011100: data = 6'b111111;
12'b1111101011101: data = 6'b111111;
12'b1111101011110: data = 6'b111111;
12'b1111101011111: data = 6'b111111;
12'b1111101100000: data = 6'b111111;
12'b1111101100001: data = 6'b101010;
12'b1111101100010: data = 6'b101010;
12'b1111101100011: data = 6'b101010;
12'b1111101100100: data = 6'b111110;
12'b1111101100101: data = 6'b111111;
12'b1111101100110: data = 6'b111110;
12'b1111101100111: data = 6'b111110;
12'b1111101101000: data = 6'b111110;
12'b1111101101001: data = 6'b111111;
12'b1111101101010: data = 6'b111111;
12'b1111101101011: data = 6'b111111;
12'b1111101101100: data = 6'b111111;
12'b1111101101101: data = 6'b111111;
12'b1111101101110: data = 6'b111111;
12'b1111101101111: data = 6'b111111;
12'b1111101110000: data = 6'b111111;
12'b1111101110001: data = 6'b111111;
12'b1111101110010: data = 6'b111111;
12'b1111101110011: data = 6'b111111;
12'b1111101110100: data = 6'b111111;
12'b1111101110101: data = 6'b111111;
12'b1111101110110: data = 6'b111111;
12'b1111101110111: data = 6'b111111;
12'b1111101111000: data = 6'b111111;
12'b1111101111001: data = 6'b111111;
12'b1111101111010: data = 6'b111111;
12'b1111101111011: data = 6'b111111;
12'b1111101111100: data = 6'b111111;
12'b1111101111101: data = 6'b111111;
12'b1111101111110: data = 6'b111111;
12'b1111101111111: data = 6'b111111;
12'b11111010000000: data = 6'b111111;
12'b11111010000001: data = 6'b111111;
12'b11111010000010: data = 6'b111111;
12'b11111010000011: data = 6'b111111;
12'b11111010000100: data = 6'b111110;
12'b11111010000101: data = 6'b111110;
12'b11111010000110: data = 6'b111110;
12'b11111010000111: data = 6'b111110;
12'b11111010001000: data = 6'b101010;
12'b11111010001001: data = 6'b010101;
12'b11111010001010: data = 6'b010101;
12'b11111010001011: data = 6'b010101;
12'b11111010001100: data = 6'b000000;
12'b11111010001101: data = 6'b000000;
12'b11111010001110: data = 6'b101010;
12'b11111010001111: data = 6'b101010;
12'b11111010010000: data = 6'b101010;
12'b11111010010001: data = 6'b101010;
12'b11111010010010: data = 6'b010101;
12'b11111010010011: data = 6'b010101;
12'b11111010010100: data = 6'b010101;
12'b11111010010101: data = 6'b010101;
12'b11111010010110: data = 6'b010101;
12'b11111010010111: data = 6'b010101;
12'b11111010011000: data = 6'b010101;
12'b11111010011001: data = 6'b010101;
12'b11111010011010: data = 6'b010101;
12'b11111010011011: data = 6'b010101;
12'b11111010011100: data = 6'b010101;
12'b11111010011101: data = 6'b010101;
12'b11111010011110: data = 6'b010101;
12'b11111010011111: data = 6'b010101;
12'b11111010100000: data = 6'b010101;
12'b11111010100001: data = 6'b010101;
12'b11111010100010: data = 6'b010101;
12'b11111010100011: data = 6'b010101;
12'b11111010100100: data = 6'b010101;
12'b11111010100101: data = 6'b010101;
12'b11111010100110: data = 6'b010101;
12'b11111010100111: data = 6'b010101;
12'b11111010101000: data = 6'b010101;
12'b11111010101001: data = 6'b010101;
12'b11111010101010: data = 6'b010101;
12'b111111000000: data = 6'b010101;
12'b111111000001: data = 6'b010101;
12'b111111000010: data = 6'b010101;
12'b111111000011: data = 6'b010101;
12'b111111000100: data = 6'b010101;
12'b111111000101: data = 6'b010101;
12'b111111000110: data = 6'b010101;
12'b111111000111: data = 6'b010101;
12'b111111001000: data = 6'b010101;
12'b111111001001: data = 6'b010101;
12'b111111001010: data = 6'b010101;
12'b111111001011: data = 6'b010101;
12'b111111001100: data = 6'b010101;
12'b111111001101: data = 6'b010101;
12'b111111001110: data = 6'b010101;
12'b111111001111: data = 6'b010101;
12'b111111010000: data = 6'b010101;
12'b111111010001: data = 6'b010101;
12'b111111010010: data = 6'b010101;
12'b111111010011: data = 6'b010101;
12'b111111010100: data = 6'b010101;
12'b111111010101: data = 6'b010101;
12'b111111010110: data = 6'b010101;
12'b111111010111: data = 6'b010101;
12'b111111011000: data = 6'b010101;
12'b111111011001: data = 6'b101010;
12'b111111011010: data = 6'b101010;
12'b111111011011: data = 6'b101010;
12'b111111011100: data = 6'b010101;
12'b111111011101: data = 6'b000000;
12'b111111011110: data = 6'b000000;
12'b111111011111: data = 6'b010101;
12'b111111100000: data = 6'b010101;
12'b111111100001: data = 6'b010101;
12'b111111100010: data = 6'b101010;
12'b111111100011: data = 6'b101010;
12'b111111100100: data = 6'b101010;
12'b111111100101: data = 6'b111110;
12'b111111100110: data = 6'b111110;
12'b111111100111: data = 6'b111111;
12'b111111101000: data = 6'b111111;
12'b111111101001: data = 6'b111111;
12'b111111101010: data = 6'b111111;
12'b111111101011: data = 6'b111111;
12'b111111101100: data = 6'b111111;
12'b111111101101: data = 6'b111111;
12'b111111101110: data = 6'b111111;
12'b111111101111: data = 6'b111111;
12'b111111110000: data = 6'b111111;
12'b111111110001: data = 6'b111111;
12'b111111110010: data = 6'b111111;
12'b111111110011: data = 6'b111111;
12'b111111110100: data = 6'b111111;
12'b111111110101: data = 6'b111111;
12'b111111110110: data = 6'b111111;
12'b111111110111: data = 6'b111111;
12'b111111111000: data = 6'b111111;
12'b111111111001: data = 6'b111111;
12'b111111111010: data = 6'b111111;
12'b111111111011: data = 6'b111111;
12'b111111111100: data = 6'b111111;
12'b111111111101: data = 6'b111111;
12'b111111111110: data = 6'b111111;
12'b111111111111: data = 6'b111111;
12'b1111111000000: data = 6'b111111;
12'b1111111000001: data = 6'b111110;
12'b1111111000010: data = 6'b101010;
12'b1111111000011: data = 6'b101010;
12'b1111111000100: data = 6'b111010;
12'b1111111000101: data = 6'b111111;
12'b1111111000110: data = 6'b111110;
12'b1111111000111: data = 6'b101010;
12'b1111111001000: data = 6'b101010;
12'b1111111001001: data = 6'b101010;
12'b1111111001010: data = 6'b111111;
12'b1111111001011: data = 6'b111111;
12'b1111111001100: data = 6'b111111;
12'b1111111001101: data = 6'b111111;
12'b1111111001110: data = 6'b111111;
12'b1111111001111: data = 6'b111111;
12'b1111111010000: data = 6'b111111;
12'b1111111010001: data = 6'b111111;
12'b1111111010010: data = 6'b111111;
12'b1111111010011: data = 6'b111111;
12'b1111111010100: data = 6'b111111;
12'b1111111010101: data = 6'b111111;
12'b1111111010110: data = 6'b111111;
12'b1111111010111: data = 6'b111111;
12'b1111111011000: data = 6'b111111;
12'b1111111011001: data = 6'b111111;
12'b1111111011010: data = 6'b111111;
12'b1111111011011: data = 6'b111111;
12'b1111111011100: data = 6'b111111;
12'b1111111011101: data = 6'b111111;
12'b1111111011110: data = 6'b111111;
12'b1111111011111: data = 6'b111111;
12'b1111111100000: data = 6'b111111;
12'b1111111100001: data = 6'b101010;
12'b1111111100010: data = 6'b101010;
12'b1111111100011: data = 6'b101010;
12'b1111111100100: data = 6'b111110;
12'b1111111100101: data = 6'b111111;
12'b1111111100110: data = 6'b111110;
12'b1111111100111: data = 6'b111110;
12'b1111111101000: data = 6'b111110;
12'b1111111101001: data = 6'b111111;
12'b1111111101010: data = 6'b111111;
12'b1111111101011: data = 6'b111111;
12'b1111111101100: data = 6'b111111;
12'b1111111101101: data = 6'b111111;
12'b1111111101110: data = 6'b111111;
12'b1111111101111: data = 6'b111111;
12'b1111111110000: data = 6'b111111;
12'b1111111110001: data = 6'b111111;
12'b1111111110010: data = 6'b111111;
12'b1111111110011: data = 6'b111111;
12'b1111111110100: data = 6'b111111;
12'b1111111110101: data = 6'b111111;
12'b1111111110110: data = 6'b111111;
12'b1111111110111: data = 6'b111111;
12'b1111111111000: data = 6'b111111;
12'b1111111111001: data = 6'b111111;
12'b1111111111010: data = 6'b111111;
12'b1111111111011: data = 6'b111111;
12'b1111111111100: data = 6'b111111;
12'b1111111111101: data = 6'b111111;
12'b1111111111110: data = 6'b111111;
12'b1111111111111: data = 6'b111111;
12'b11111110000000: data = 6'b111111;
12'b11111110000001: data = 6'b111111;
12'b11111110000010: data = 6'b111111;
12'b11111110000011: data = 6'b111111;
12'b11111110000100: data = 6'b111110;
12'b11111110000101: data = 6'b111110;
12'b11111110000110: data = 6'b111110;
12'b11111110000111: data = 6'b111110;
12'b11111110001000: data = 6'b101010;
12'b11111110001001: data = 6'b010101;
12'b11111110001010: data = 6'b010101;
12'b11111110001011: data = 6'b010101;
12'b11111110001100: data = 6'b000000;
12'b11111110001101: data = 6'b000000;
12'b11111110001110: data = 6'b101010;
12'b11111110001111: data = 6'b101010;
12'b11111110010000: data = 6'b101010;
12'b11111110010001: data = 6'b101010;
12'b11111110010010: data = 6'b010101;
12'b11111110010011: data = 6'b010101;
12'b11111110010100: data = 6'b010101;
12'b11111110010101: data = 6'b010101;
12'b11111110010110: data = 6'b010101;
12'b11111110010111: data = 6'b010101;
12'b11111110011000: data = 6'b010101;
12'b11111110011001: data = 6'b010101;
12'b11111110011010: data = 6'b010101;
12'b11111110011011: data = 6'b010101;
12'b11111110011100: data = 6'b010101;
12'b11111110011101: data = 6'b010101;
12'b11111110011110: data = 6'b010101;
12'b11111110011111: data = 6'b010101;
12'b11111110100000: data = 6'b010101;
12'b11111110100001: data = 6'b010101;
12'b11111110100010: data = 6'b010101;
12'b11111110100011: data = 6'b010101;
12'b11111110100100: data = 6'b010101;
12'b11111110100101: data = 6'b010101;
12'b11111110100110: data = 6'b010101;
12'b11111110100111: data = 6'b010101;
12'b11111110101000: data = 6'b010101;
12'b11111110101001: data = 6'b010101;
12'b11111110101010: data = 6'b010101;
12'b1000000000000: data = 6'b010101;
12'b1000000000001: data = 6'b010101;
12'b1000000000010: data = 6'b010101;
12'b1000000000011: data = 6'b010101;
12'b1000000000100: data = 6'b010101;
12'b1000000000101: data = 6'b010101;
12'b1000000000110: data = 6'b010101;
12'b1000000000111: data = 6'b010101;
12'b1000000001000: data = 6'b010101;
12'b1000000001001: data = 6'b010101;
12'b1000000001010: data = 6'b010101;
12'b1000000001011: data = 6'b010101;
12'b1000000001100: data = 6'b010101;
12'b1000000001101: data = 6'b010101;
12'b1000000001110: data = 6'b010101;
12'b1000000001111: data = 6'b010101;
12'b1000000010000: data = 6'b010101;
12'b1000000010001: data = 6'b010101;
12'b1000000010010: data = 6'b010101;
12'b1000000010011: data = 6'b010101;
12'b1000000010100: data = 6'b010101;
12'b1000000010101: data = 6'b010101;
12'b1000000010110: data = 6'b010101;
12'b1000000010111: data = 6'b010101;
12'b1000000011000: data = 6'b010101;
12'b1000000011001: data = 6'b101010;
12'b1000000011010: data = 6'b101010;
12'b1000000011011: data = 6'b101010;
12'b1000000011100: data = 6'b010101;
12'b1000000011101: data = 6'b000000;
12'b1000000011110: data = 6'b000000;
12'b1000000011111: data = 6'b010101;
12'b1000000100000: data = 6'b010101;
12'b1000000100001: data = 6'b010101;
12'b1000000100010: data = 6'b101010;
12'b1000000100011: data = 6'b111010;
12'b1000000100100: data = 6'b111010;
12'b1000000100101: data = 6'b111111;
12'b1000000100110: data = 6'b111110;
12'b1000000100111: data = 6'b111111;
12'b1000000101000: data = 6'b111111;
12'b1000000101001: data = 6'b111111;
12'b1000000101010: data = 6'b111111;
12'b1000000101011: data = 6'b111111;
12'b1000000101100: data = 6'b111111;
12'b1000000101101: data = 6'b111111;
12'b1000000101110: data = 6'b111111;
12'b1000000101111: data = 6'b111111;
12'b1000000110000: data = 6'b111111;
12'b1000000110001: data = 6'b111111;
12'b1000000110010: data = 6'b111111;
12'b1000000110011: data = 6'b111111;
12'b1000000110100: data = 6'b111111;
12'b1000000110101: data = 6'b111111;
12'b1000000110110: data = 6'b111111;
12'b1000000110111: data = 6'b111111;
12'b1000000111000: data = 6'b111111;
12'b1000000111001: data = 6'b111111;
12'b1000000111010: data = 6'b111111;
12'b1000000111011: data = 6'b111111;
12'b1000000111100: data = 6'b111111;
12'b1000000111101: data = 6'b111111;
12'b1000000111110: data = 6'b111111;
12'b1000000111111: data = 6'b111111;
12'b10000001000000: data = 6'b111111;
12'b10000001000001: data = 6'b111111;
12'b10000001000010: data = 6'b111110;
12'b10000001000011: data = 6'b111010;
12'b10000001000100: data = 6'b111110;
12'b10000001000101: data = 6'b111110;
12'b10000001000110: data = 6'b111110;
12'b10000001000111: data = 6'b101010;
12'b10000001001000: data = 6'b101010;
12'b10000001001001: data = 6'b101010;
12'b10000001001010: data = 6'b111111;
12'b10000001001011: data = 6'b111111;
12'b10000001001100: data = 6'b111111;
12'b10000001001101: data = 6'b111111;
12'b10000001001110: data = 6'b111111;
12'b10000001001111: data = 6'b111111;
12'b10000001010000: data = 6'b111111;
12'b10000001010001: data = 6'b111111;
12'b10000001010010: data = 6'b111111;
12'b10000001010011: data = 6'b111111;
12'b10000001010100: data = 6'b111111;
12'b10000001010101: data = 6'b111111;
12'b10000001010110: data = 6'b111111;
12'b10000001010111: data = 6'b111111;
12'b10000001011000: data = 6'b111111;
12'b10000001011001: data = 6'b111111;
12'b10000001011010: data = 6'b111111;
12'b10000001011011: data = 6'b111111;
12'b10000001011100: data = 6'b111111;
12'b10000001011101: data = 6'b111111;
12'b10000001011110: data = 6'b111111;
12'b10000001011111: data = 6'b111111;
12'b10000001100000: data = 6'b111111;
12'b10000001100001: data = 6'b101010;
12'b10000001100010: data = 6'b101010;
12'b10000001100011: data = 6'b101010;
12'b10000001100100: data = 6'b111111;
12'b10000001100101: data = 6'b111111;
12'b10000001100110: data = 6'b111111;
12'b10000001100111: data = 6'b111110;
12'b10000001101000: data = 6'b111111;
12'b10000001101001: data = 6'b111111;
12'b10000001101010: data = 6'b111111;
12'b10000001101011: data = 6'b111111;
12'b10000001101100: data = 6'b111111;
12'b10000001101101: data = 6'b111111;
12'b10000001101110: data = 6'b111111;
12'b10000001101111: data = 6'b111111;
12'b10000001110000: data = 6'b111111;
12'b10000001110001: data = 6'b111111;
12'b10000001110010: data = 6'b111111;
12'b10000001110011: data = 6'b111111;
12'b10000001110100: data = 6'b111111;
12'b10000001110101: data = 6'b111111;
12'b10000001110110: data = 6'b111111;
12'b10000001110111: data = 6'b111111;
12'b10000001111000: data = 6'b111111;
12'b10000001111001: data = 6'b111111;
12'b10000001111010: data = 6'b111111;
12'b10000001111011: data = 6'b111111;
12'b10000001111100: data = 6'b111111;
12'b10000001111101: data = 6'b111111;
12'b10000001111110: data = 6'b111111;
12'b10000001111111: data = 6'b111111;
12'b100000010000000: data = 6'b111111;
12'b100000010000001: data = 6'b111111;
12'b100000010000010: data = 6'b111111;
12'b100000010000011: data = 6'b111111;
12'b100000010000100: data = 6'b111111;
12'b100000010000101: data = 6'b111111;
12'b100000010000110: data = 6'b111110;
12'b100000010000111: data = 6'b111010;
12'b100000010001000: data = 6'b101010;
12'b100000010001001: data = 6'b010101;
12'b100000010001010: data = 6'b010101;
12'b100000010001011: data = 6'b010101;
12'b100000010001100: data = 6'b000000;
12'b100000010001101: data = 6'b000000;
12'b100000010001110: data = 6'b101010;
12'b100000010001111: data = 6'b101010;
12'b100000010010000: data = 6'b101010;
12'b100000010010001: data = 6'b101010;
12'b100000010010010: data = 6'b010101;
12'b100000010010011: data = 6'b010101;
12'b100000010010100: data = 6'b010101;
12'b100000010010101: data = 6'b010101;
12'b100000010010110: data = 6'b010101;
12'b100000010010111: data = 6'b010101;
12'b100000010011000: data = 6'b010101;
12'b100000010011001: data = 6'b010101;
12'b100000010011010: data = 6'b010101;
12'b100000010011011: data = 6'b010101;
12'b100000010011100: data = 6'b010101;
12'b100000010011101: data = 6'b010101;
12'b100000010011110: data = 6'b010101;
12'b100000010011111: data = 6'b010101;
12'b100000010100000: data = 6'b010101;
12'b100000010100001: data = 6'b010101;
12'b100000010100010: data = 6'b010101;
12'b100000010100011: data = 6'b010101;
12'b100000010100100: data = 6'b010101;
12'b100000010100101: data = 6'b010101;
12'b100000010100110: data = 6'b010101;
12'b100000010100111: data = 6'b010101;
12'b100000010101000: data = 6'b010101;
12'b100000010101001: data = 6'b010101;
12'b100000010101010: data = 6'b010101;
12'b1000001000000: data = 6'b010101;
12'b1000001000001: data = 6'b010101;
12'b1000001000010: data = 6'b010101;
12'b1000001000011: data = 6'b010101;
12'b1000001000100: data = 6'b010101;
12'b1000001000101: data = 6'b010101;
12'b1000001000110: data = 6'b010101;
12'b1000001000111: data = 6'b010101;
12'b1000001001000: data = 6'b010101;
12'b1000001001001: data = 6'b010101;
12'b1000001001010: data = 6'b010101;
12'b1000001001011: data = 6'b010101;
12'b1000001001100: data = 6'b010101;
12'b1000001001101: data = 6'b010101;
12'b1000001001110: data = 6'b010101;
12'b1000001001111: data = 6'b010101;
12'b1000001010000: data = 6'b010101;
12'b1000001010001: data = 6'b010101;
12'b1000001010010: data = 6'b010101;
12'b1000001010011: data = 6'b010101;
12'b1000001010100: data = 6'b010101;
12'b1000001010101: data = 6'b010101;
12'b1000001010110: data = 6'b010101;
12'b1000001010111: data = 6'b010101;
12'b1000001011000: data = 6'b010101;
12'b1000001011001: data = 6'b101010;
12'b1000001011010: data = 6'b101010;
12'b1000001011011: data = 6'b101010;
12'b1000001011100: data = 6'b010101;
12'b1000001011101: data = 6'b000000;
12'b1000001011110: data = 6'b000000;
12'b1000001011111: data = 6'b010101;
12'b1000001100000: data = 6'b010101;
12'b1000001100001: data = 6'b010101;
12'b1000001100010: data = 6'b101010;
12'b1000001100011: data = 6'b111110;
12'b1000001100100: data = 6'b111110;
12'b1000001100101: data = 6'b111111;
12'b1000001100110: data = 6'b111111;
12'b1000001100111: data = 6'b111111;
12'b1000001101000: data = 6'b111111;
12'b1000001101001: data = 6'b111111;
12'b1000001101010: data = 6'b111111;
12'b1000001101011: data = 6'b111111;
12'b1000001101100: data = 6'b111111;
12'b1000001101101: data = 6'b111111;
12'b1000001101110: data = 6'b111111;
12'b1000001101111: data = 6'b111111;
12'b1000001110000: data = 6'b111111;
12'b1000001110001: data = 6'b111111;
12'b1000001110010: data = 6'b111111;
12'b1000001110011: data = 6'b111111;
12'b1000001110100: data = 6'b111111;
12'b1000001110101: data = 6'b111111;
12'b1000001110110: data = 6'b111111;
12'b1000001110111: data = 6'b111111;
12'b1000001111000: data = 6'b111111;
12'b1000001111001: data = 6'b111111;
12'b1000001111010: data = 6'b111111;
12'b1000001111011: data = 6'b111111;
12'b1000001111100: data = 6'b111111;
12'b1000001111101: data = 6'b111111;
12'b1000001111110: data = 6'b111111;
12'b1000001111111: data = 6'b111111;
12'b10000011000000: data = 6'b111111;
12'b10000011000001: data = 6'b111111;
12'b10000011000010: data = 6'b111110;
12'b10000011000011: data = 6'b111110;
12'b10000011000100: data = 6'b111110;
12'b10000011000101: data = 6'b101010;
12'b10000011000110: data = 6'b101010;
12'b10000011000111: data = 6'b101010;
12'b10000011001000: data = 6'b101010;
12'b10000011001001: data = 6'b101010;
12'b10000011001010: data = 6'b111111;
12'b10000011001011: data = 6'b111111;
12'b10000011001100: data = 6'b111111;
12'b10000011001101: data = 6'b111111;
12'b10000011001110: data = 6'b111111;
12'b10000011001111: data = 6'b111111;
12'b10000011010000: data = 6'b111111;
12'b10000011010001: data = 6'b111111;
12'b10000011010010: data = 6'b111111;
12'b10000011010011: data = 6'b111111;
12'b10000011010100: data = 6'b111111;
12'b10000011010101: data = 6'b111111;
12'b10000011010110: data = 6'b111111;
12'b10000011010111: data = 6'b111111;
12'b10000011011000: data = 6'b111111;
12'b10000011011001: data = 6'b111111;
12'b10000011011010: data = 6'b111111;
12'b10000011011011: data = 6'b111111;
12'b10000011011100: data = 6'b111111;
12'b10000011011101: data = 6'b111111;
12'b10000011011110: data = 6'b111111;
12'b10000011011111: data = 6'b111111;
12'b10000011100000: data = 6'b111111;
12'b10000011100001: data = 6'b101010;
12'b10000011100010: data = 6'b101010;
12'b10000011100011: data = 6'b101010;
12'b10000011100100: data = 6'b111111;
12'b10000011100101: data = 6'b111111;
12'b10000011100110: data = 6'b111111;
12'b10000011100111: data = 6'b111111;
12'b10000011101000: data = 6'b111111;
12'b10000011101001: data = 6'b111111;
12'b10000011101010: data = 6'b111111;
12'b10000011101011: data = 6'b111111;
12'b10000011101100: data = 6'b111111;
12'b10000011101101: data = 6'b111111;
12'b10000011101110: data = 6'b111111;
12'b10000011101111: data = 6'b111111;
12'b10000011110000: data = 6'b111111;
12'b10000011110001: data = 6'b111111;
12'b10000011110010: data = 6'b111111;
12'b10000011110011: data = 6'b111111;
12'b10000011110100: data = 6'b111111;
12'b10000011110101: data = 6'b111111;
12'b10000011110110: data = 6'b111111;
12'b10000011110111: data = 6'b111111;
12'b10000011111000: data = 6'b111111;
12'b10000011111001: data = 6'b111111;
12'b10000011111010: data = 6'b111111;
12'b10000011111011: data = 6'b111111;
12'b10000011111100: data = 6'b111111;
12'b10000011111101: data = 6'b111111;
12'b10000011111110: data = 6'b111111;
12'b10000011111111: data = 6'b111111;
12'b100000110000000: data = 6'b111111;
12'b100000110000001: data = 6'b111111;
12'b100000110000010: data = 6'b111111;
12'b100000110000011: data = 6'b111111;
12'b100000110000100: data = 6'b111111;
12'b100000110000101: data = 6'b111111;
12'b100000110000110: data = 6'b101010;
12'b100000110000111: data = 6'b111010;
12'b100000110001000: data = 6'b101010;
12'b100000110001001: data = 6'b010101;
12'b100000110001010: data = 6'b010101;
12'b100000110001011: data = 6'b010101;
12'b100000110001100: data = 6'b000000;
12'b100000110001101: data = 6'b000000;
12'b100000110001110: data = 6'b101010;
12'b100000110001111: data = 6'b101010;
12'b100000110010000: data = 6'b101010;
12'b100000110010001: data = 6'b101010;
12'b100000110010010: data = 6'b010101;
12'b100000110010011: data = 6'b010101;
12'b100000110010100: data = 6'b010101;
12'b100000110010101: data = 6'b010101;
12'b100000110010110: data = 6'b010101;
12'b100000110010111: data = 6'b010101;
12'b100000110011000: data = 6'b010101;
12'b100000110011001: data = 6'b010101;
12'b100000110011010: data = 6'b010101;
12'b100000110011011: data = 6'b010101;
12'b100000110011100: data = 6'b010101;
12'b100000110011101: data = 6'b010101;
12'b100000110011110: data = 6'b010101;
12'b100000110011111: data = 6'b010101;
12'b100000110100000: data = 6'b010101;
12'b100000110100001: data = 6'b010101;
12'b100000110100010: data = 6'b010101;
12'b100000110100011: data = 6'b010101;
12'b100000110100100: data = 6'b010101;
12'b100000110100101: data = 6'b010101;
12'b100000110100110: data = 6'b010101;
12'b100000110100111: data = 6'b010101;
12'b100000110101000: data = 6'b010101;
12'b100000110101001: data = 6'b010101;
12'b100000110101010: data = 6'b010101;
12'b1000010000000: data = 6'b010101;
12'b1000010000001: data = 6'b010101;
12'b1000010000010: data = 6'b010101;
12'b1000010000011: data = 6'b010101;
12'b1000010000100: data = 6'b010101;
12'b1000010000101: data = 6'b010101;
12'b1000010000110: data = 6'b010101;
12'b1000010000111: data = 6'b010101;
12'b1000010001000: data = 6'b010101;
12'b1000010001001: data = 6'b010101;
12'b1000010001010: data = 6'b010101;
12'b1000010001011: data = 6'b010101;
12'b1000010001100: data = 6'b010101;
12'b1000010001101: data = 6'b010101;
12'b1000010001110: data = 6'b010101;
12'b1000010001111: data = 6'b010101;
12'b1000010010000: data = 6'b010101;
12'b1000010010001: data = 6'b010101;
12'b1000010010010: data = 6'b010101;
12'b1000010010011: data = 6'b010101;
12'b1000010010100: data = 6'b010101;
12'b1000010010101: data = 6'b010101;
12'b1000010010110: data = 6'b010101;
12'b1000010010111: data = 6'b010101;
12'b1000010011000: data = 6'b010101;
12'b1000010011001: data = 6'b101010;
12'b1000010011010: data = 6'b101010;
12'b1000010011011: data = 6'b101010;
12'b1000010011100: data = 6'b010101;
12'b1000010011101: data = 6'b000000;
12'b1000010011110: data = 6'b000000;
12'b1000010011111: data = 6'b010101;
12'b1000010100000: data = 6'b010101;
12'b1000010100001: data = 6'b010101;
12'b1000010100010: data = 6'b101010;
12'b1000010100011: data = 6'b111110;
12'b1000010100100: data = 6'b101010;
12'b1000010100101: data = 6'b111111;
12'b1000010100110: data = 6'b111111;
12'b1000010100111: data = 6'b111111;
12'b1000010101000: data = 6'b111111;
12'b1000010101001: data = 6'b111111;
12'b1000010101010: data = 6'b111111;
12'b1000010101011: data = 6'b111111;
12'b1000010101100: data = 6'b111111;
12'b1000010101101: data = 6'b111111;
12'b1000010101110: data = 6'b111111;
12'b1000010101111: data = 6'b111111;
12'b1000010110000: data = 6'b111111;
12'b1000010110001: data = 6'b111111;
12'b1000010110010: data = 6'b111111;
12'b1000010110011: data = 6'b111111;
12'b1000010110100: data = 6'b111111;
12'b1000010110101: data = 6'b111111;
12'b1000010110110: data = 6'b111111;
12'b1000010110111: data = 6'b111111;
12'b1000010111000: data = 6'b111111;
12'b1000010111001: data = 6'b111111;
12'b1000010111010: data = 6'b111111;
12'b1000010111011: data = 6'b111111;
12'b1000010111100: data = 6'b111111;
12'b1000010111101: data = 6'b111111;
12'b1000010111110: data = 6'b111111;
12'b1000010111111: data = 6'b111111;
12'b10000101000000: data = 6'b111111;
12'b10000101000001: data = 6'b111111;
12'b10000101000010: data = 6'b111110;
12'b10000101000011: data = 6'b111111;
12'b10000101000100: data = 6'b111110;
12'b10000101000101: data = 6'b111111;
12'b10000101000110: data = 6'b101010;
12'b10000101000111: data = 6'b101010;
12'b10000101001000: data = 6'b101010;
12'b10000101001001: data = 6'b101010;
12'b10000101001010: data = 6'b111111;
12'b10000101001011: data = 6'b111111;
12'b10000101001100: data = 6'b111111;
12'b10000101001101: data = 6'b111111;
12'b10000101001110: data = 6'b111111;
12'b10000101001111: data = 6'b111111;
12'b10000101010000: data = 6'b111111;
12'b10000101010001: data = 6'b111111;
12'b10000101010010: data = 6'b111111;
12'b10000101010011: data = 6'b111111;
12'b10000101010100: data = 6'b111111;
12'b10000101010101: data = 6'b111111;
12'b10000101010110: data = 6'b111111;
12'b10000101010111: data = 6'b111111;
12'b10000101011000: data = 6'b111111;
12'b10000101011001: data = 6'b111111;
12'b10000101011010: data = 6'b111111;
12'b10000101011011: data = 6'b111111;
12'b10000101011100: data = 6'b111111;
12'b10000101011101: data = 6'b111111;
12'b10000101011110: data = 6'b111111;
12'b10000101011111: data = 6'b111111;
12'b10000101100000: data = 6'b111111;
12'b10000101100001: data = 6'b101010;
12'b10000101100010: data = 6'b101010;
12'b10000101100011: data = 6'b101010;
12'b10000101100100: data = 6'b111111;
12'b10000101100101: data = 6'b111111;
12'b10000101100110: data = 6'b111111;
12'b10000101100111: data = 6'b111111;
12'b10000101101000: data = 6'b111111;
12'b10000101101001: data = 6'b111111;
12'b10000101101010: data = 6'b111111;
12'b10000101101011: data = 6'b111111;
12'b10000101101100: data = 6'b111111;
12'b10000101101101: data = 6'b111111;
12'b10000101101110: data = 6'b111111;
12'b10000101101111: data = 6'b111111;
12'b10000101110000: data = 6'b111111;
12'b10000101110001: data = 6'b111111;
12'b10000101110010: data = 6'b111111;
12'b10000101110011: data = 6'b111111;
12'b10000101110100: data = 6'b111111;
12'b10000101110101: data = 6'b111111;
12'b10000101110110: data = 6'b111111;
12'b10000101110111: data = 6'b111111;
12'b10000101111000: data = 6'b111111;
12'b10000101111001: data = 6'b111111;
12'b10000101111010: data = 6'b111111;
12'b10000101111011: data = 6'b111111;
12'b10000101111100: data = 6'b111111;
12'b10000101111101: data = 6'b111111;
12'b10000101111110: data = 6'b111111;
12'b10000101111111: data = 6'b111111;
12'b100001010000000: data = 6'b111111;
12'b100001010000001: data = 6'b111111;
12'b100001010000010: data = 6'b111111;
12'b100001010000011: data = 6'b111111;
12'b100001010000100: data = 6'b111111;
12'b100001010000101: data = 6'b111111;
12'b100001010000110: data = 6'b101010;
12'b100001010000111: data = 6'b101010;
12'b100001010001000: data = 6'b101010;
12'b100001010001001: data = 6'b010101;
12'b100001010001010: data = 6'b010101;
12'b100001010001011: data = 6'b010101;
12'b100001010001100: data = 6'b000000;
12'b100001010001101: data = 6'b000000;
12'b100001010001110: data = 6'b101010;
12'b100001010001111: data = 6'b101010;
12'b100001010010000: data = 6'b101010;
12'b100001010010001: data = 6'b101010;
12'b100001010010010: data = 6'b010101;
12'b100001010010011: data = 6'b010101;
12'b100001010010100: data = 6'b010101;
12'b100001010010101: data = 6'b010101;
12'b100001010010110: data = 6'b010101;
12'b100001010010111: data = 6'b010101;
12'b100001010011000: data = 6'b010101;
12'b100001010011001: data = 6'b010101;
12'b100001010011010: data = 6'b010101;
12'b100001010011011: data = 6'b010101;
12'b100001010011100: data = 6'b010101;
12'b100001010011101: data = 6'b010101;
12'b100001010011110: data = 6'b010101;
12'b100001010011111: data = 6'b010101;
12'b100001010100000: data = 6'b010101;
12'b100001010100001: data = 6'b010101;
12'b100001010100010: data = 6'b010101;
12'b100001010100011: data = 6'b010101;
12'b100001010100100: data = 6'b010101;
12'b100001010100101: data = 6'b010101;
12'b100001010100110: data = 6'b010101;
12'b100001010100111: data = 6'b010101;
12'b100001010101000: data = 6'b010101;
12'b100001010101001: data = 6'b010101;
12'b100001010101010: data = 6'b010101;
12'b1000011000000: data = 6'b010101;
12'b1000011000001: data = 6'b010101;
12'b1000011000010: data = 6'b010101;
12'b1000011000011: data = 6'b010101;
12'b1000011000100: data = 6'b010101;
12'b1000011000101: data = 6'b010101;
12'b1000011000110: data = 6'b010101;
12'b1000011000111: data = 6'b010101;
12'b1000011001000: data = 6'b010101;
12'b1000011001001: data = 6'b010101;
12'b1000011001010: data = 6'b010101;
12'b1000011001011: data = 6'b010101;
12'b1000011001100: data = 6'b010101;
12'b1000011001101: data = 6'b010101;
12'b1000011001110: data = 6'b010101;
12'b1000011001111: data = 6'b010101;
12'b1000011010000: data = 6'b010101;
12'b1000011010001: data = 6'b010101;
12'b1000011010010: data = 6'b010101;
12'b1000011010011: data = 6'b010101;
12'b1000011010100: data = 6'b010101;
12'b1000011010101: data = 6'b010101;
12'b1000011010110: data = 6'b010101;
12'b1000011010111: data = 6'b010101;
12'b1000011011000: data = 6'b010101;
12'b1000011011001: data = 6'b101010;
12'b1000011011010: data = 6'b101010;
12'b1000011011011: data = 6'b101010;
12'b1000011011100: data = 6'b010101;
12'b1000011011101: data = 6'b000000;
12'b1000011011110: data = 6'b000000;
12'b1000011011111: data = 6'b010101;
12'b1000011100000: data = 6'b010101;
12'b1000011100001: data = 6'b010101;
12'b1000011100010: data = 6'b101010;
12'b1000011100011: data = 6'b101010;
12'b1000011100100: data = 6'b101010;
12'b1000011100101: data = 6'b111111;
12'b1000011100110: data = 6'b111111;
12'b1000011100111: data = 6'b111111;
12'b1000011101000: data = 6'b111111;
12'b1000011101001: data = 6'b111111;
12'b1000011101010: data = 6'b111111;
12'b1000011101011: data = 6'b111111;
12'b1000011101100: data = 6'b111111;
12'b1000011101101: data = 6'b111111;
12'b1000011101110: data = 6'b111111;
12'b1000011101111: data = 6'b111111;
12'b1000011110000: data = 6'b111111;
12'b1000011110001: data = 6'b111111;
12'b1000011110010: data = 6'b111111;
12'b1000011110011: data = 6'b111111;
12'b1000011110100: data = 6'b111111;
12'b1000011110101: data = 6'b111111;
12'b1000011110110: data = 6'b111111;
12'b1000011110111: data = 6'b111111;
12'b1000011111000: data = 6'b111111;
12'b1000011111001: data = 6'b111111;
12'b1000011111010: data = 6'b111111;
12'b1000011111011: data = 6'b111111;
12'b1000011111100: data = 6'b111111;
12'b1000011111101: data = 6'b111111;
12'b1000011111110: data = 6'b111111;
12'b1000011111111: data = 6'b111111;
12'b10000111000000: data = 6'b111111;
12'b10000111000001: data = 6'b111111;
12'b10000111000010: data = 6'b111111;
12'b10000111000011: data = 6'b101010;
12'b10000111000100: data = 6'b111111;
12'b10000111000101: data = 6'b111111;
12'b10000111000110: data = 6'b101010;
12'b10000111000111: data = 6'b101010;
12'b10000111001000: data = 6'b101010;
12'b10000111001001: data = 6'b101010;
12'b10000111001010: data = 6'b111111;
12'b10000111001011: data = 6'b111111;
12'b10000111001100: data = 6'b111111;
12'b10000111001101: data = 6'b111111;
12'b10000111001110: data = 6'b111111;
12'b10000111001111: data = 6'b111111;
12'b10000111010000: data = 6'b111111;
12'b10000111010001: data = 6'b111111;
12'b10000111010010: data = 6'b111111;
12'b10000111010011: data = 6'b111111;
12'b10000111010100: data = 6'b111111;
12'b10000111010101: data = 6'b111111;
12'b10000111010110: data = 6'b111111;
12'b10000111010111: data = 6'b111111;
12'b10000111011000: data = 6'b111111;
12'b10000111011001: data = 6'b111111;
12'b10000111011010: data = 6'b111111;
12'b10000111011011: data = 6'b111111;
12'b10000111011100: data = 6'b111111;
12'b10000111011101: data = 6'b111111;
12'b10000111011110: data = 6'b111111;
12'b10000111011111: data = 6'b111111;
12'b10000111100000: data = 6'b111111;
12'b10000111100001: data = 6'b101010;
12'b10000111100010: data = 6'b101010;
12'b10000111100011: data = 6'b101010;
12'b10000111100100: data = 6'b101010;
12'b10000111100101: data = 6'b111111;
12'b10000111100110: data = 6'b111111;
12'b10000111100111: data = 6'b111111;
12'b10000111101000: data = 6'b111111;
12'b10000111101001: data = 6'b111111;
12'b10000111101010: data = 6'b111111;
12'b10000111101011: data = 6'b111111;
12'b10000111101100: data = 6'b111111;
12'b10000111101101: data = 6'b111111;
12'b10000111101110: data = 6'b111111;
12'b10000111101111: data = 6'b111111;
12'b10000111110000: data = 6'b111111;
12'b10000111110001: data = 6'b111111;
12'b10000111110010: data = 6'b111111;
12'b10000111110011: data = 6'b111111;
12'b10000111110100: data = 6'b111111;
12'b10000111110101: data = 6'b111111;
12'b10000111110110: data = 6'b111111;
12'b10000111110111: data = 6'b111111;
12'b10000111111000: data = 6'b111111;
12'b10000111111001: data = 6'b111111;
12'b10000111111010: data = 6'b111111;
12'b10000111111011: data = 6'b111111;
12'b10000111111100: data = 6'b111111;
12'b10000111111101: data = 6'b111111;
12'b10000111111110: data = 6'b111111;
12'b10000111111111: data = 6'b111111;
12'b100001110000000: data = 6'b111111;
12'b100001110000001: data = 6'b111111;
12'b100001110000010: data = 6'b111111;
12'b100001110000011: data = 6'b111111;
12'b100001110000100: data = 6'b111111;
12'b100001110000101: data = 6'b111111;
12'b100001110000110: data = 6'b101010;
12'b100001110000111: data = 6'b101010;
12'b100001110001000: data = 6'b101010;
12'b100001110001001: data = 6'b010101;
12'b100001110001010: data = 6'b010101;
12'b100001110001011: data = 6'b010101;
12'b100001110001100: data = 6'b000000;
12'b100001110001101: data = 6'b000000;
12'b100001110001110: data = 6'b101010;
12'b100001110001111: data = 6'b101010;
12'b100001110010000: data = 6'b101010;
12'b100001110010001: data = 6'b101010;
12'b100001110010010: data = 6'b010101;
12'b100001110010011: data = 6'b010101;
12'b100001110010100: data = 6'b010101;
12'b100001110010101: data = 6'b010101;
12'b100001110010110: data = 6'b010101;
12'b100001110010111: data = 6'b010101;
12'b100001110011000: data = 6'b010101;
12'b100001110011001: data = 6'b010101;
12'b100001110011010: data = 6'b010101;
12'b100001110011011: data = 6'b010101;
12'b100001110011100: data = 6'b010101;
12'b100001110011101: data = 6'b010101;
12'b100001110011110: data = 6'b010101;
12'b100001110011111: data = 6'b010101;
12'b100001110100000: data = 6'b010101;
12'b100001110100001: data = 6'b010101;
12'b100001110100010: data = 6'b010101;
12'b100001110100011: data = 6'b010101;
12'b100001110100100: data = 6'b010101;
12'b100001110100101: data = 6'b010101;
12'b100001110100110: data = 6'b010101;
12'b100001110100111: data = 6'b010101;
12'b100001110101000: data = 6'b010101;
12'b100001110101001: data = 6'b010101;
12'b100001110101010: data = 6'b010101;
12'b1000100000000: data = 6'b010101;
12'b1000100000001: data = 6'b010101;
12'b1000100000010: data = 6'b010101;
12'b1000100000011: data = 6'b010101;
12'b1000100000100: data = 6'b010101;
12'b1000100000101: data = 6'b010101;
12'b1000100000110: data = 6'b010101;
12'b1000100000111: data = 6'b010101;
12'b1000100001000: data = 6'b010101;
12'b1000100001001: data = 6'b010101;
12'b1000100001010: data = 6'b010101;
12'b1000100001011: data = 6'b010101;
12'b1000100001100: data = 6'b010101;
12'b1000100001101: data = 6'b010101;
12'b1000100001110: data = 6'b010101;
12'b1000100001111: data = 6'b010101;
12'b1000100010000: data = 6'b010101;
12'b1000100010001: data = 6'b010101;
12'b1000100010010: data = 6'b010101;
12'b1000100010011: data = 6'b010101;
12'b1000100010100: data = 6'b010101;
12'b1000100010101: data = 6'b010101;
12'b1000100010110: data = 6'b010101;
12'b1000100010111: data = 6'b010101;
12'b1000100011000: data = 6'b010101;
12'b1000100011001: data = 6'b101010;
12'b1000100011010: data = 6'b101010;
12'b1000100011011: data = 6'b101010;
12'b1000100011100: data = 6'b010101;
12'b1000100011101: data = 6'b000000;
12'b1000100011110: data = 6'b000000;
12'b1000100011111: data = 6'b010101;
12'b1000100100000: data = 6'b010101;
12'b1000100100001: data = 6'b010101;
12'b1000100100010: data = 6'b101010;
12'b1000100100011: data = 6'b101010;
12'b1000100100100: data = 6'b101010;
12'b1000100100101: data = 6'b111111;
12'b1000100100110: data = 6'b111111;
12'b1000100100111: data = 6'b111111;
12'b1000100101000: data = 6'b111111;
12'b1000100101001: data = 6'b111111;
12'b1000100101010: data = 6'b111111;
12'b1000100101011: data = 6'b111111;
12'b1000100101100: data = 6'b111111;
12'b1000100101101: data = 6'b111111;
12'b1000100101110: data = 6'b111111;
12'b1000100101111: data = 6'b111111;
12'b1000100110000: data = 6'b111111;
12'b1000100110001: data = 6'b111111;
12'b1000100110010: data = 6'b111111;
12'b1000100110011: data = 6'b111111;
12'b1000100110100: data = 6'b111111;
12'b1000100110101: data = 6'b111111;
12'b1000100110110: data = 6'b111111;
12'b1000100110111: data = 6'b111111;
12'b1000100111000: data = 6'b111111;
12'b1000100111001: data = 6'b111111;
12'b1000100111010: data = 6'b111111;
12'b1000100111011: data = 6'b111111;
12'b1000100111100: data = 6'b111111;
12'b1000100111101: data = 6'b111111;
12'b1000100111110: data = 6'b111111;
12'b1000100111111: data = 6'b111111;
12'b10001001000000: data = 6'b111111;
12'b10001001000001: data = 6'b111111;
12'b10001001000010: data = 6'b111111;
12'b10001001000011: data = 6'b111111;
12'b10001001000100: data = 6'b111111;
12'b10001001000101: data = 6'b111111;
12'b10001001000110: data = 6'b101010;
12'b10001001000111: data = 6'b101010;
12'b10001001001000: data = 6'b101010;
12'b10001001001001: data = 6'b101010;
12'b10001001001010: data = 6'b111111;
12'b10001001001011: data = 6'b111111;
12'b10001001001100: data = 6'b111111;
12'b10001001001101: data = 6'b111111;
12'b10001001001110: data = 6'b111111;
12'b10001001001111: data = 6'b111111;
12'b10001001010000: data = 6'b111111;
12'b10001001010001: data = 6'b111111;
12'b10001001010010: data = 6'b111111;
12'b10001001010011: data = 6'b111111;
12'b10001001010100: data = 6'b111111;
12'b10001001010101: data = 6'b111111;
12'b10001001010110: data = 6'b111111;
12'b10001001010111: data = 6'b111111;
12'b10001001011000: data = 6'b111111;
12'b10001001011001: data = 6'b111111;
12'b10001001011010: data = 6'b111111;
12'b10001001011011: data = 6'b111111;
12'b10001001011100: data = 6'b111111;
12'b10001001011101: data = 6'b111111;
12'b10001001011110: data = 6'b111111;
12'b10001001011111: data = 6'b111111;
12'b10001001100000: data = 6'b111111;
12'b10001001100001: data = 6'b101010;
12'b10001001100010: data = 6'b101010;
12'b10001001100011: data = 6'b101010;
12'b10001001100100: data = 6'b101010;
12'b10001001100101: data = 6'b111111;
12'b10001001100110: data = 6'b111111;
12'b10001001100111: data = 6'b111111;
12'b10001001101000: data = 6'b111111;
12'b10001001101001: data = 6'b111111;
12'b10001001101010: data = 6'b111111;
12'b10001001101011: data = 6'b111111;
12'b10001001101100: data = 6'b111111;
12'b10001001101101: data = 6'b111111;
12'b10001001101110: data = 6'b111111;
12'b10001001101111: data = 6'b111111;
12'b10001001110000: data = 6'b111111;
12'b10001001110001: data = 6'b111111;
12'b10001001110010: data = 6'b111111;
12'b10001001110011: data = 6'b111111;
12'b10001001110100: data = 6'b111111;
12'b10001001110101: data = 6'b111111;
12'b10001001110110: data = 6'b111111;
12'b10001001110111: data = 6'b111111;
12'b10001001111000: data = 6'b111111;
12'b10001001111001: data = 6'b111111;
12'b10001001111010: data = 6'b111111;
12'b10001001111011: data = 6'b111111;
12'b10001001111100: data = 6'b111111;
12'b10001001111101: data = 6'b111111;
12'b10001001111110: data = 6'b111111;
12'b10001001111111: data = 6'b111111;
12'b100010010000000: data = 6'b111111;
12'b100010010000001: data = 6'b111111;
12'b100010010000010: data = 6'b111111;
12'b100010010000011: data = 6'b111111;
12'b100010010000100: data = 6'b111111;
12'b100010010000101: data = 6'b101010;
12'b100010010000110: data = 6'b101010;
12'b100010010000111: data = 6'b101010;
12'b100010010001000: data = 6'b101010;
12'b100010010001001: data = 6'b010101;
12'b100010010001010: data = 6'b010101;
12'b100010010001011: data = 6'b010101;
12'b100010010001100: data = 6'b000000;
12'b100010010001101: data = 6'b000000;
12'b100010010001110: data = 6'b101010;
12'b100010010001111: data = 6'b101010;
12'b100010010010000: data = 6'b101010;
12'b100010010010001: data = 6'b101010;
12'b100010010010010: data = 6'b010101;
12'b100010010010011: data = 6'b010101;
12'b100010010010100: data = 6'b010101;
12'b100010010010101: data = 6'b010101;
12'b100010010010110: data = 6'b010101;
12'b100010010010111: data = 6'b010101;
12'b100010010011000: data = 6'b010101;
12'b100010010011001: data = 6'b010101;
12'b100010010011010: data = 6'b010101;
12'b100010010011011: data = 6'b010101;
12'b100010010011100: data = 6'b010101;
12'b100010010011101: data = 6'b010101;
12'b100010010011110: data = 6'b010101;
12'b100010010011111: data = 6'b010101;
12'b100010010100000: data = 6'b010101;
12'b100010010100001: data = 6'b010101;
12'b100010010100010: data = 6'b010101;
12'b100010010100011: data = 6'b010101;
12'b100010010100100: data = 6'b010101;
12'b100010010100101: data = 6'b010101;
12'b100010010100110: data = 6'b010101;
12'b100010010100111: data = 6'b010101;
12'b100010010101000: data = 6'b010101;
12'b100010010101001: data = 6'b010101;
12'b100010010101010: data = 6'b010101;
12'b1000101000000: data = 6'b010101;
12'b1000101000001: data = 6'b010101;
12'b1000101000010: data = 6'b010101;
12'b1000101000011: data = 6'b010101;
12'b1000101000100: data = 6'b010101;
12'b1000101000101: data = 6'b010101;
12'b1000101000110: data = 6'b010101;
12'b1000101000111: data = 6'b010101;
12'b1000101001000: data = 6'b010101;
12'b1000101001001: data = 6'b010101;
12'b1000101001010: data = 6'b010101;
12'b1000101001011: data = 6'b010101;
12'b1000101001100: data = 6'b010101;
12'b1000101001101: data = 6'b010101;
12'b1000101001110: data = 6'b010101;
12'b1000101001111: data = 6'b010101;
12'b1000101010000: data = 6'b010101;
12'b1000101010001: data = 6'b010101;
12'b1000101010010: data = 6'b010101;
12'b1000101010011: data = 6'b010101;
12'b1000101010100: data = 6'b010101;
12'b1000101010101: data = 6'b010101;
12'b1000101010110: data = 6'b010101;
12'b1000101010111: data = 6'b010101;
12'b1000101011000: data = 6'b010101;
12'b1000101011001: data = 6'b101010;
12'b1000101011010: data = 6'b101010;
12'b1000101011011: data = 6'b101010;
12'b1000101011100: data = 6'b010101;
12'b1000101011101: data = 6'b000000;
12'b1000101011110: data = 6'b000000;
12'b1000101011111: data = 6'b010101;
12'b1000101100000: data = 6'b010101;
12'b1000101100001: data = 6'b010101;
12'b1000101100010: data = 6'b101010;
12'b1000101100011: data = 6'b101010;
12'b1000101100100: data = 6'b101010;
12'b1000101100101: data = 6'b101010;
12'b1000101100110: data = 6'b101010;
12'b1000101100111: data = 6'b111111;
12'b1000101101000: data = 6'b111111;
12'b1000101101001: data = 6'b111111;
12'b1000101101010: data = 6'b111111;
12'b1000101101011: data = 6'b111111;
12'b1000101101100: data = 6'b111111;
12'b1000101101101: data = 6'b111111;
12'b1000101101110: data = 6'b111111;
12'b1000101101111: data = 6'b111111;
12'b1000101110000: data = 6'b111111;
12'b1000101110001: data = 6'b111111;
12'b1000101110010: data = 6'b111111;
12'b1000101110011: data = 6'b111111;
12'b1000101110100: data = 6'b111111;
12'b1000101110101: data = 6'b111111;
12'b1000101110110: data = 6'b111111;
12'b1000101110111: data = 6'b111111;
12'b1000101111000: data = 6'b111111;
12'b1000101111001: data = 6'b111111;
12'b1000101111010: data = 6'b111111;
12'b1000101111011: data = 6'b111111;
12'b1000101111100: data = 6'b111111;
12'b1000101111101: data = 6'b111111;
12'b1000101111110: data = 6'b111111;
12'b1000101111111: data = 6'b111111;
12'b10001011000000: data = 6'b111111;
12'b10001011000001: data = 6'b111111;
12'b10001011000010: data = 6'b101010;
12'b10001011000011: data = 6'b101010;
12'b10001011000100: data = 6'b101010;
12'b10001011000101: data = 6'b101010;
12'b10001011000110: data = 6'b101010;
12'b10001011000111: data = 6'b101010;
12'b10001011001000: data = 6'b101010;
12'b10001011001001: data = 6'b101010;
12'b10001011001010: data = 6'b111111;
12'b10001011001011: data = 6'b111111;
12'b10001011001100: data = 6'b111111;
12'b10001011001101: data = 6'b111111;
12'b10001011001110: data = 6'b111111;
12'b10001011001111: data = 6'b111111;
12'b10001011010000: data = 6'b111111;
12'b10001011010001: data = 6'b111111;
12'b10001011010010: data = 6'b111111;
12'b10001011010011: data = 6'b111111;
12'b10001011010100: data = 6'b111111;
12'b10001011010101: data = 6'b111111;
12'b10001011010110: data = 6'b111111;
12'b10001011010111: data = 6'b111111;
12'b10001011011000: data = 6'b111111;
12'b10001011011001: data = 6'b111111;
12'b10001011011010: data = 6'b111111;
12'b10001011011011: data = 6'b111111;
12'b10001011011100: data = 6'b111111;
12'b10001011011101: data = 6'b111111;
12'b10001011011110: data = 6'b111111;
12'b10001011011111: data = 6'b111111;
12'b10001011100000: data = 6'b111111;
12'b10001011100001: data = 6'b101010;
12'b10001011100010: data = 6'b101010;
12'b10001011100011: data = 6'b101010;
12'b10001011100100: data = 6'b101010;
12'b10001011100101: data = 6'b101010;
12'b10001011100110: data = 6'b101010;
12'b10001011100111: data = 6'b101010;
12'b10001011101000: data = 6'b101010;
12'b10001011101001: data = 6'b111111;
12'b10001011101010: data = 6'b111111;
12'b10001011101011: data = 6'b111111;
12'b10001011101100: data = 6'b111111;
12'b10001011101101: data = 6'b111111;
12'b10001011101110: data = 6'b111111;
12'b10001011101111: data = 6'b111111;
12'b10001011110000: data = 6'b111111;
12'b10001011110001: data = 6'b111111;
12'b10001011110010: data = 6'b111111;
12'b10001011110011: data = 6'b111111;
12'b10001011110100: data = 6'b111111;
12'b10001011110101: data = 6'b111111;
12'b10001011110110: data = 6'b111111;
12'b10001011110111: data = 6'b111111;
12'b10001011111000: data = 6'b111111;
12'b10001011111001: data = 6'b111111;
12'b10001011111010: data = 6'b111111;
12'b10001011111011: data = 6'b111111;
12'b10001011111100: data = 6'b111111;
12'b10001011111101: data = 6'b111111;
12'b10001011111110: data = 6'b111111;
12'b10001011111111: data = 6'b111111;
12'b100010110000000: data = 6'b111111;
12'b100010110000001: data = 6'b111111;
12'b100010110000010: data = 6'b111111;
12'b100010110000011: data = 6'b111111;
12'b100010110000100: data = 6'b101010;
12'b100010110000101: data = 6'b101010;
12'b100010110000110: data = 6'b101010;
12'b100010110000111: data = 6'b101010;
12'b100010110001000: data = 6'b101010;
12'b100010110001001: data = 6'b010101;
12'b100010110001010: data = 6'b010101;
12'b100010110001011: data = 6'b010101;
12'b100010110001100: data = 6'b000000;
12'b100010110001101: data = 6'b000000;
12'b100010110001110: data = 6'b101010;
12'b100010110001111: data = 6'b101010;
12'b100010110010000: data = 6'b101010;
12'b100010110010001: data = 6'b101010;
12'b100010110010010: data = 6'b010101;
12'b100010110010011: data = 6'b010101;
12'b100010110010100: data = 6'b010101;
12'b100010110010101: data = 6'b010101;
12'b100010110010110: data = 6'b010101;
12'b100010110010111: data = 6'b010101;
12'b100010110011000: data = 6'b010101;
12'b100010110011001: data = 6'b010101;
12'b100010110011010: data = 6'b010101;
12'b100010110011011: data = 6'b010101;
12'b100010110011100: data = 6'b010101;
12'b100010110011101: data = 6'b010101;
12'b100010110011110: data = 6'b010101;
12'b100010110011111: data = 6'b010101;
12'b100010110100000: data = 6'b010101;
12'b100010110100001: data = 6'b010101;
12'b100010110100010: data = 6'b010101;
12'b100010110100011: data = 6'b010101;
12'b100010110100100: data = 6'b010101;
12'b100010110100101: data = 6'b010101;
12'b100010110100110: data = 6'b010101;
12'b100010110100111: data = 6'b010101;
12'b100010110101000: data = 6'b010101;
12'b100010110101001: data = 6'b010101;
12'b100010110101010: data = 6'b010101;
12'b1000110000000: data = 6'b010101;
12'b1000110000001: data = 6'b010101;
12'b1000110000010: data = 6'b010101;
12'b1000110000011: data = 6'b010101;
12'b1000110000100: data = 6'b010101;
12'b1000110000101: data = 6'b010101;
12'b1000110000110: data = 6'b010101;
12'b1000110000111: data = 6'b010101;
12'b1000110001000: data = 6'b010101;
12'b1000110001001: data = 6'b010101;
12'b1000110001010: data = 6'b010101;
12'b1000110001011: data = 6'b010101;
12'b1000110001100: data = 6'b010101;
12'b1000110001101: data = 6'b010101;
12'b1000110001110: data = 6'b010101;
12'b1000110001111: data = 6'b010101;
12'b1000110010000: data = 6'b010101;
12'b1000110010001: data = 6'b010101;
12'b1000110010010: data = 6'b010101;
12'b1000110010011: data = 6'b010101;
12'b1000110010100: data = 6'b010101;
12'b1000110010101: data = 6'b010101;
12'b1000110010110: data = 6'b010101;
12'b1000110010111: data = 6'b010101;
12'b1000110011000: data = 6'b010101;
12'b1000110011001: data = 6'b101010;
12'b1000110011010: data = 6'b101010;
12'b1000110011011: data = 6'b101010;
12'b1000110011100: data = 6'b010101;
12'b1000110011101: data = 6'b000000;
12'b1000110011110: data = 6'b000000;
12'b1000110011111: data = 6'b010101;
12'b1000110100000: data = 6'b010101;
12'b1000110100001: data = 6'b010101;
12'b1000110100010: data = 6'b101010;
12'b1000110100011: data = 6'b101010;
12'b1000110100100: data = 6'b101010;
12'b1000110100101: data = 6'b101010;
12'b1000110100110: data = 6'b101010;
12'b1000110100111: data = 6'b111111;
12'b1000110101000: data = 6'b111111;
12'b1000110101001: data = 6'b111111;
12'b1000110101010: data = 6'b111111;
12'b1000110101011: data = 6'b111111;
12'b1000110101100: data = 6'b111111;
12'b1000110101101: data = 6'b111111;
12'b1000110101110: data = 6'b111111;
12'b1000110101111: data = 6'b111111;
12'b1000110110000: data = 6'b111111;
12'b1000110110001: data = 6'b111111;
12'b1000110110010: data = 6'b111111;
12'b1000110110011: data = 6'b111111;
12'b1000110110100: data = 6'b111111;
12'b1000110110101: data = 6'b111111;
12'b1000110110110: data = 6'b111111;
12'b1000110110111: data = 6'b111111;
12'b1000110111000: data = 6'b111111;
12'b1000110111001: data = 6'b111111;
12'b1000110111010: data = 6'b111111;
12'b1000110111011: data = 6'b111111;
12'b1000110111100: data = 6'b111111;
12'b1000110111101: data = 6'b111111;
12'b1000110111110: data = 6'b111111;
12'b1000110111111: data = 6'b111111;
12'b10001101000000: data = 6'b111111;
12'b10001101000001: data = 6'b111111;
12'b10001101000010: data = 6'b101010;
12'b10001101000011: data = 6'b101010;
12'b10001101000100: data = 6'b101010;
12'b10001101000101: data = 6'b101010;
12'b10001101000110: data = 6'b101010;
12'b10001101000111: data = 6'b101010;
12'b10001101001000: data = 6'b101010;
12'b10001101001001: data = 6'b101010;
12'b10001101001010: data = 6'b111111;
12'b10001101001011: data = 6'b111111;
12'b10001101001100: data = 6'b111111;
12'b10001101001101: data = 6'b111111;
12'b10001101001110: data = 6'b111111;
12'b10001101001111: data = 6'b111111;
12'b10001101010000: data = 6'b111111;
12'b10001101010001: data = 6'b111111;
12'b10001101010010: data = 6'b111111;
12'b10001101010011: data = 6'b111111;
12'b10001101010100: data = 6'b111111;
12'b10001101010101: data = 6'b111111;
12'b10001101010110: data = 6'b111111;
12'b10001101010111: data = 6'b111111;
12'b10001101011000: data = 6'b111111;
12'b10001101011001: data = 6'b111111;
12'b10001101011010: data = 6'b111111;
12'b10001101011011: data = 6'b111111;
12'b10001101011100: data = 6'b111111;
12'b10001101011101: data = 6'b111111;
12'b10001101011110: data = 6'b111111;
12'b10001101011111: data = 6'b111111;
12'b10001101100000: data = 6'b111111;
12'b10001101100001: data = 6'b101010;
12'b10001101100010: data = 6'b101010;
12'b10001101100011: data = 6'b101010;
12'b10001101100100: data = 6'b101010;
12'b10001101100101: data = 6'b101010;
12'b10001101100110: data = 6'b101010;
12'b10001101100111: data = 6'b101010;
12'b10001101101000: data = 6'b101010;
12'b10001101101001: data = 6'b111111;
12'b10001101101010: data = 6'b111111;
12'b10001101101011: data = 6'b111111;
12'b10001101101100: data = 6'b111111;
12'b10001101101101: data = 6'b111111;
12'b10001101101110: data = 6'b111111;
12'b10001101101111: data = 6'b111111;
12'b10001101110000: data = 6'b111111;
12'b10001101110001: data = 6'b111111;
12'b10001101110010: data = 6'b111111;
12'b10001101110011: data = 6'b111111;
12'b10001101110100: data = 6'b111111;
12'b10001101110101: data = 6'b111111;
12'b10001101110110: data = 6'b111111;
12'b10001101110111: data = 6'b111111;
12'b10001101111000: data = 6'b111111;
12'b10001101111001: data = 6'b111111;
12'b10001101111010: data = 6'b111111;
12'b10001101111011: data = 6'b111111;
12'b10001101111100: data = 6'b111111;
12'b10001101111101: data = 6'b111111;
12'b10001101111110: data = 6'b111111;
12'b10001101111111: data = 6'b111111;
12'b100011010000000: data = 6'b111111;
12'b100011010000001: data = 6'b111111;
12'b100011010000010: data = 6'b111111;
12'b100011010000011: data = 6'b111111;
12'b100011010000100: data = 6'b101010;
12'b100011010000101: data = 6'b101010;
12'b100011010000110: data = 6'b101010;
12'b100011010000111: data = 6'b101010;
12'b100011010001000: data = 6'b101010;
12'b100011010001001: data = 6'b010101;
12'b100011010001010: data = 6'b010101;
12'b100011010001011: data = 6'b010101;
12'b100011010001100: data = 6'b000000;
12'b100011010001101: data = 6'b000000;
12'b100011010001110: data = 6'b101010;
12'b100011010001111: data = 6'b101010;
12'b100011010010000: data = 6'b101010;
12'b100011010010001: data = 6'b101010;
12'b100011010010010: data = 6'b010101;
12'b100011010010011: data = 6'b010101;
12'b100011010010100: data = 6'b010101;
12'b100011010010101: data = 6'b010101;
12'b100011010010110: data = 6'b010101;
12'b100011010010111: data = 6'b010101;
12'b100011010011000: data = 6'b010101;
12'b100011010011001: data = 6'b010101;
12'b100011010011010: data = 6'b010101;
12'b100011010011011: data = 6'b010101;
12'b100011010011100: data = 6'b010101;
12'b100011010011101: data = 6'b010101;
12'b100011010011110: data = 6'b010101;
12'b100011010011111: data = 6'b010101;
12'b100011010100000: data = 6'b010101;
12'b100011010100001: data = 6'b010101;
12'b100011010100010: data = 6'b010101;
12'b100011010100011: data = 6'b010101;
12'b100011010100100: data = 6'b010101;
12'b100011010100101: data = 6'b010101;
12'b100011010100110: data = 6'b010101;
12'b100011010100111: data = 6'b010101;
12'b100011010101000: data = 6'b010101;
12'b100011010101001: data = 6'b010101;
12'b100011010101010: data = 6'b010101;
12'b1000111000000: data = 6'b010101;
12'b1000111000001: data = 6'b010101;
12'b1000111000010: data = 6'b010101;
12'b1000111000011: data = 6'b010101;
12'b1000111000100: data = 6'b010101;
12'b1000111000101: data = 6'b010101;
12'b1000111000110: data = 6'b010101;
12'b1000111000111: data = 6'b010101;
12'b1000111001000: data = 6'b010101;
12'b1000111001001: data = 6'b010101;
12'b1000111001010: data = 6'b010101;
12'b1000111001011: data = 6'b010101;
12'b1000111001100: data = 6'b010101;
12'b1000111001101: data = 6'b010101;
12'b1000111001110: data = 6'b010101;
12'b1000111001111: data = 6'b010101;
12'b1000111010000: data = 6'b010101;
12'b1000111010001: data = 6'b010101;
12'b1000111010010: data = 6'b010101;
12'b1000111010011: data = 6'b010101;
12'b1000111010100: data = 6'b010101;
12'b1000111010101: data = 6'b010101;
12'b1000111010110: data = 6'b010101;
12'b1000111010111: data = 6'b010101;
12'b1000111011000: data = 6'b010101;
12'b1000111011001: data = 6'b101010;
12'b1000111011010: data = 6'b101010;
12'b1000111011011: data = 6'b101010;
12'b1000111011100: data = 6'b010101;
12'b1000111011101: data = 6'b000000;
12'b1000111011110: data = 6'b000000;
12'b1000111011111: data = 6'b010101;
12'b1000111100000: data = 6'b010101;
12'b1000111100001: data = 6'b010101;
12'b1000111100010: data = 6'b101010;
12'b1000111100011: data = 6'b101010;
12'b1000111100100: data = 6'b101010;
12'b1000111100101: data = 6'b101010;
12'b1000111100110: data = 6'b101010;
12'b1000111100111: data = 6'b111111;
12'b1000111101000: data = 6'b111111;
12'b1000111101001: data = 6'b111111;
12'b1000111101010: data = 6'b111111;
12'b1000111101011: data = 6'b111111;
12'b1000111101100: data = 6'b111111;
12'b1000111101101: data = 6'b111111;
12'b1000111101110: data = 6'b111111;
12'b1000111101111: data = 6'b111111;
12'b1000111110000: data = 6'b111111;
12'b1000111110001: data = 6'b111111;
12'b1000111110010: data = 6'b111111;
12'b1000111110011: data = 6'b111111;
12'b1000111110100: data = 6'b111111;
12'b1000111110101: data = 6'b111111;
12'b1000111110110: data = 6'b111111;
12'b1000111110111: data = 6'b111111;
12'b1000111111000: data = 6'b111111;
12'b1000111111001: data = 6'b111111;
12'b1000111111010: data = 6'b111111;
12'b1000111111011: data = 6'b111111;
12'b1000111111100: data = 6'b111111;
12'b1000111111101: data = 6'b111111;
12'b1000111111110: data = 6'b111111;
12'b1000111111111: data = 6'b111111;
12'b10001111000000: data = 6'b111111;
12'b10001111000001: data = 6'b111111;
12'b10001111000010: data = 6'b101010;
12'b10001111000011: data = 6'b101010;
12'b10001111000100: data = 6'b101010;
12'b10001111000101: data = 6'b101010;
12'b10001111000110: data = 6'b101010;
12'b10001111000111: data = 6'b101010;
12'b10001111001000: data = 6'b101010;
12'b10001111001001: data = 6'b101010;
12'b10001111001010: data = 6'b111111;
12'b10001111001011: data = 6'b111111;
12'b10001111001100: data = 6'b111111;
12'b10001111001101: data = 6'b111111;
12'b10001111001110: data = 6'b111111;
12'b10001111001111: data = 6'b111111;
12'b10001111010000: data = 6'b111111;
12'b10001111010001: data = 6'b111111;
12'b10001111010010: data = 6'b111111;
12'b10001111010011: data = 6'b111111;
12'b10001111010100: data = 6'b111111;
12'b10001111010101: data = 6'b111111;
12'b10001111010110: data = 6'b111111;
12'b10001111010111: data = 6'b111111;
12'b10001111011000: data = 6'b111111;
12'b10001111011001: data = 6'b111111;
12'b10001111011010: data = 6'b111111;
12'b10001111011011: data = 6'b111111;
12'b10001111011100: data = 6'b111111;
12'b10001111011101: data = 6'b111111;
12'b10001111011110: data = 6'b111111;
12'b10001111011111: data = 6'b111111;
12'b10001111100000: data = 6'b111111;
12'b10001111100001: data = 6'b101010;
12'b10001111100010: data = 6'b101010;
12'b10001111100011: data = 6'b101010;
12'b10001111100100: data = 6'b101010;
12'b10001111100101: data = 6'b101010;
12'b10001111100110: data = 6'b101010;
12'b10001111100111: data = 6'b101010;
12'b10001111101000: data = 6'b101010;
12'b10001111101001: data = 6'b111111;
12'b10001111101010: data = 6'b111111;
12'b10001111101011: data = 6'b111111;
12'b10001111101100: data = 6'b111111;
12'b10001111101101: data = 6'b111111;
12'b10001111101110: data = 6'b111111;
12'b10001111101111: data = 6'b111111;
12'b10001111110000: data = 6'b111111;
12'b10001111110001: data = 6'b111111;
12'b10001111110010: data = 6'b111111;
12'b10001111110011: data = 6'b111111;
12'b10001111110100: data = 6'b111111;
12'b10001111110101: data = 6'b111111;
12'b10001111110110: data = 6'b111111;
12'b10001111110111: data = 6'b111111;
12'b10001111111000: data = 6'b111111;
12'b10001111111001: data = 6'b111111;
12'b10001111111010: data = 6'b111111;
12'b10001111111011: data = 6'b111111;
12'b10001111111100: data = 6'b111111;
12'b10001111111101: data = 6'b111111;
12'b10001111111110: data = 6'b111111;
12'b10001111111111: data = 6'b111111;
12'b100011110000000: data = 6'b111111;
12'b100011110000001: data = 6'b111111;
12'b100011110000010: data = 6'b111111;
12'b100011110000011: data = 6'b111111;
12'b100011110000100: data = 6'b101010;
12'b100011110000101: data = 6'b101010;
12'b100011110000110: data = 6'b101010;
12'b100011110000111: data = 6'b101010;
12'b100011110001000: data = 6'b101010;
12'b100011110001001: data = 6'b010101;
12'b100011110001010: data = 6'b010101;
12'b100011110001011: data = 6'b010101;
12'b100011110001100: data = 6'b000000;
12'b100011110001101: data = 6'b000000;
12'b100011110001110: data = 6'b101010;
12'b100011110001111: data = 6'b101010;
12'b100011110010000: data = 6'b101010;
12'b100011110010001: data = 6'b101010;
12'b100011110010010: data = 6'b010101;
12'b100011110010011: data = 6'b010101;
12'b100011110010100: data = 6'b010101;
12'b100011110010101: data = 6'b010101;
12'b100011110010110: data = 6'b010101;
12'b100011110010111: data = 6'b010101;
12'b100011110011000: data = 6'b010101;
12'b100011110011001: data = 6'b010101;
12'b100011110011010: data = 6'b010101;
12'b100011110011011: data = 6'b010101;
12'b100011110011100: data = 6'b010101;
12'b100011110011101: data = 6'b010101;
12'b100011110011110: data = 6'b010101;
12'b100011110011111: data = 6'b010101;
12'b100011110100000: data = 6'b010101;
12'b100011110100001: data = 6'b010101;
12'b100011110100010: data = 6'b010101;
12'b100011110100011: data = 6'b010101;
12'b100011110100100: data = 6'b010101;
12'b100011110100101: data = 6'b010101;
12'b100011110100110: data = 6'b010101;
12'b100011110100111: data = 6'b010101;
12'b100011110101000: data = 6'b010101;
12'b100011110101001: data = 6'b010101;
12'b100011110101010: data = 6'b010101;
12'b1001000000000: data = 6'b010101;
12'b1001000000001: data = 6'b010101;
12'b1001000000010: data = 6'b010101;
12'b1001000000011: data = 6'b010101;
12'b1001000000100: data = 6'b010101;
12'b1001000000101: data = 6'b010101;
12'b1001000000110: data = 6'b010101;
12'b1001000000111: data = 6'b010101;
12'b1001000001000: data = 6'b010101;
12'b1001000001001: data = 6'b010101;
12'b1001000001010: data = 6'b010101;
12'b1001000001011: data = 6'b010101;
12'b1001000001100: data = 6'b010101;
12'b1001000001101: data = 6'b010101;
12'b1001000001110: data = 6'b010101;
12'b1001000001111: data = 6'b010101;
12'b1001000010000: data = 6'b010101;
12'b1001000010001: data = 6'b010101;
12'b1001000010010: data = 6'b010101;
12'b1001000010011: data = 6'b010101;
12'b1001000010100: data = 6'b010101;
12'b1001000010101: data = 6'b010101;
12'b1001000010110: data = 6'b010101;
12'b1001000010111: data = 6'b010101;
12'b1001000011000: data = 6'b010101;
12'b1001000011001: data = 6'b101010;
12'b1001000011010: data = 6'b101010;
12'b1001000011011: data = 6'b101010;
12'b1001000011100: data = 6'b010101;
12'b1001000011101: data = 6'b000000;
12'b1001000011110: data = 6'b000000;
12'b1001000011111: data = 6'b010101;
12'b1001000100000: data = 6'b010101;
12'b1001000100001: data = 6'b010101;
12'b1001000100010: data = 6'b101010;
12'b1001000100011: data = 6'b101010;
12'b1001000100100: data = 6'b101010;
12'b1001000100101: data = 6'b101010;
12'b1001000100110: data = 6'b101010;
12'b1001000100111: data = 6'b111111;
12'b1001000101000: data = 6'b111111;
12'b1001000101001: data = 6'b111111;
12'b1001000101010: data = 6'b111111;
12'b1001000101011: data = 6'b111111;
12'b1001000101100: data = 6'b111111;
12'b1001000101101: data = 6'b111111;
12'b1001000101110: data = 6'b111111;
12'b1001000101111: data = 6'b111111;
12'b1001000110000: data = 6'b111111;
12'b1001000110001: data = 6'b111111;
12'b1001000110010: data = 6'b111111;
12'b1001000110011: data = 6'b111111;
12'b1001000110100: data = 6'b111111;
12'b1001000110101: data = 6'b111111;
12'b1001000110110: data = 6'b111111;
12'b1001000110111: data = 6'b111111;
12'b1001000111000: data = 6'b111111;
12'b1001000111001: data = 6'b111111;
12'b1001000111010: data = 6'b111111;
12'b1001000111011: data = 6'b111111;
12'b1001000111100: data = 6'b111111;
12'b1001000111101: data = 6'b111111;
12'b1001000111110: data = 6'b111111;
12'b1001000111111: data = 6'b111111;
12'b10010001000000: data = 6'b111111;
12'b10010001000001: data = 6'b111111;
12'b10010001000010: data = 6'b101010;
12'b10010001000011: data = 6'b101010;
12'b10010001000100: data = 6'b101010;
12'b10010001000101: data = 6'b101010;
12'b10010001000110: data = 6'b101010;
12'b10010001000111: data = 6'b101010;
12'b10010001001000: data = 6'b101010;
12'b10010001001001: data = 6'b101010;
12'b10010001001010: data = 6'b111111;
12'b10010001001011: data = 6'b111111;
12'b10010001001100: data = 6'b111111;
12'b10010001001101: data = 6'b111111;
12'b10010001001110: data = 6'b111111;
12'b10010001001111: data = 6'b111111;
12'b10010001010000: data = 6'b111111;
12'b10010001010001: data = 6'b111111;
12'b10010001010010: data = 6'b111111;
12'b10010001010011: data = 6'b111111;
12'b10010001010100: data = 6'b111111;
12'b10010001010101: data = 6'b111111;
12'b10010001010110: data = 6'b111111;
12'b10010001010111: data = 6'b111111;
12'b10010001011000: data = 6'b111111;
12'b10010001011001: data = 6'b111111;
12'b10010001011010: data = 6'b111111;
12'b10010001011011: data = 6'b111111;
12'b10010001011100: data = 6'b111111;
12'b10010001011101: data = 6'b111111;
12'b10010001011110: data = 6'b111111;
12'b10010001011111: data = 6'b111111;
12'b10010001100000: data = 6'b111111;
12'b10010001100001: data = 6'b101010;
12'b10010001100010: data = 6'b101010;
12'b10010001100011: data = 6'b101010;
12'b10010001100100: data = 6'b101010;
12'b10010001100101: data = 6'b101010;
12'b10010001100110: data = 6'b101010;
12'b10010001100111: data = 6'b101010;
12'b10010001101000: data = 6'b101010;
12'b10010001101001: data = 6'b111111;
12'b10010001101010: data = 6'b111111;
12'b10010001101011: data = 6'b111111;
12'b10010001101100: data = 6'b111111;
12'b10010001101101: data = 6'b111111;
12'b10010001101110: data = 6'b111111;
12'b10010001101111: data = 6'b111111;
12'b10010001110000: data = 6'b111111;
12'b10010001110001: data = 6'b111111;
12'b10010001110010: data = 6'b111111;
12'b10010001110011: data = 6'b111111;
12'b10010001110100: data = 6'b111111;
12'b10010001110101: data = 6'b111111;
12'b10010001110110: data = 6'b111111;
12'b10010001110111: data = 6'b111111;
12'b10010001111000: data = 6'b111111;
12'b10010001111001: data = 6'b111111;
12'b10010001111010: data = 6'b111111;
12'b10010001111011: data = 6'b111111;
12'b10010001111100: data = 6'b111111;
12'b10010001111101: data = 6'b111111;
12'b10010001111110: data = 6'b111111;
12'b10010001111111: data = 6'b111111;
12'b100100010000000: data = 6'b111111;
12'b100100010000001: data = 6'b111111;
12'b100100010000010: data = 6'b111111;
12'b100100010000011: data = 6'b111111;
12'b100100010000100: data = 6'b101010;
12'b100100010000101: data = 6'b101010;
12'b100100010000110: data = 6'b101010;
12'b100100010000111: data = 6'b101010;
12'b100100010001000: data = 6'b101010;
12'b100100010001001: data = 6'b010101;
12'b100100010001010: data = 6'b010101;
12'b100100010001011: data = 6'b010101;
12'b100100010001100: data = 6'b000000;
12'b100100010001101: data = 6'b000000;
12'b100100010001110: data = 6'b101010;
12'b100100010001111: data = 6'b101010;
12'b100100010010000: data = 6'b101010;
12'b100100010010001: data = 6'b101010;
12'b100100010010010: data = 6'b010101;
12'b100100010010011: data = 6'b010101;
12'b100100010010100: data = 6'b010101;
12'b100100010010101: data = 6'b010101;
12'b100100010010110: data = 6'b010101;
12'b100100010010111: data = 6'b010101;
12'b100100010011000: data = 6'b010101;
12'b100100010011001: data = 6'b010101;
12'b100100010011010: data = 6'b010101;
12'b100100010011011: data = 6'b010101;
12'b100100010011100: data = 6'b010101;
12'b100100010011101: data = 6'b010101;
12'b100100010011110: data = 6'b010101;
12'b100100010011111: data = 6'b010101;
12'b100100010100000: data = 6'b010101;
12'b100100010100001: data = 6'b010101;
12'b100100010100010: data = 6'b010101;
12'b100100010100011: data = 6'b010101;
12'b100100010100100: data = 6'b010101;
12'b100100010100101: data = 6'b010101;
12'b100100010100110: data = 6'b010101;
12'b100100010100111: data = 6'b010101;
12'b100100010101000: data = 6'b010101;
12'b100100010101001: data = 6'b010101;
12'b100100010101010: data = 6'b010101;
12'b1001001000000: data = 6'b010101;
12'b1001001000001: data = 6'b010101;
12'b1001001000010: data = 6'b010101;
12'b1001001000011: data = 6'b010101;
12'b1001001000100: data = 6'b010101;
12'b1001001000101: data = 6'b010101;
12'b1001001000110: data = 6'b010101;
12'b1001001000111: data = 6'b010101;
12'b1001001001000: data = 6'b010101;
12'b1001001001001: data = 6'b010101;
12'b1001001001010: data = 6'b010101;
12'b1001001001011: data = 6'b010101;
12'b1001001001100: data = 6'b010101;
12'b1001001001101: data = 6'b010101;
12'b1001001001110: data = 6'b010101;
12'b1001001001111: data = 6'b010101;
12'b1001001010000: data = 6'b010101;
12'b1001001010001: data = 6'b010101;
12'b1001001010010: data = 6'b010101;
12'b1001001010011: data = 6'b010101;
12'b1001001010100: data = 6'b010101;
12'b1001001010101: data = 6'b010101;
12'b1001001010110: data = 6'b010101;
12'b1001001010111: data = 6'b010101;
12'b1001001011000: data = 6'b010101;
12'b1001001011001: data = 6'b101010;
12'b1001001011010: data = 6'b101010;
12'b1001001011011: data = 6'b101010;
12'b1001001011100: data = 6'b010101;
12'b1001001011101: data = 6'b000000;
12'b1001001011110: data = 6'b000000;
12'b1001001011111: data = 6'b010101;
12'b1001001100000: data = 6'b010101;
12'b1001001100001: data = 6'b010101;
12'b1001001100010: data = 6'b101010;
12'b1001001100011: data = 6'b101010;
12'b1001001100100: data = 6'b101010;
12'b1001001100101: data = 6'b101010;
12'b1001001100110: data = 6'b101010;
12'b1001001100111: data = 6'b111111;
12'b1001001101000: data = 6'b111111;
12'b1001001101001: data = 6'b111111;
12'b1001001101010: data = 6'b111111;
12'b1001001101011: data = 6'b111111;
12'b1001001101100: data = 6'b111111;
12'b1001001101101: data = 6'b111111;
12'b1001001101110: data = 6'b111111;
12'b1001001101111: data = 6'b111111;
12'b1001001110000: data = 6'b111111;
12'b1001001110001: data = 6'b111111;
12'b1001001110010: data = 6'b111111;
12'b1001001110011: data = 6'b111111;
12'b1001001110100: data = 6'b111111;
12'b1001001110101: data = 6'b111111;
12'b1001001110110: data = 6'b111111;
12'b1001001110111: data = 6'b111111;
12'b1001001111000: data = 6'b111111;
12'b1001001111001: data = 6'b111111;
12'b1001001111010: data = 6'b111111;
12'b1001001111011: data = 6'b111111;
12'b1001001111100: data = 6'b111111;
12'b1001001111101: data = 6'b111111;
12'b1001001111110: data = 6'b111111;
12'b1001001111111: data = 6'b111111;
12'b10010011000000: data = 6'b111111;
12'b10010011000001: data = 6'b111111;
12'b10010011000010: data = 6'b101010;
12'b10010011000011: data = 6'b101010;
12'b10010011000100: data = 6'b101010;
12'b10010011000101: data = 6'b101010;
12'b10010011000110: data = 6'b101010;
12'b10010011000111: data = 6'b101010;
12'b10010011001000: data = 6'b101010;
12'b10010011001001: data = 6'b101010;
12'b10010011001010: data = 6'b111111;
12'b10010011001011: data = 6'b111111;
12'b10010011001100: data = 6'b111111;
12'b10010011001101: data = 6'b111111;
12'b10010011001110: data = 6'b111111;
12'b10010011001111: data = 6'b111111;
12'b10010011010000: data = 6'b111111;
12'b10010011010001: data = 6'b111111;
12'b10010011010010: data = 6'b111111;
12'b10010011010011: data = 6'b111111;
12'b10010011010100: data = 6'b111111;
12'b10010011010101: data = 6'b111111;
12'b10010011010110: data = 6'b111111;
12'b10010011010111: data = 6'b111111;
12'b10010011011000: data = 6'b111111;
12'b10010011011001: data = 6'b111111;
12'b10010011011010: data = 6'b111111;
12'b10010011011011: data = 6'b111111;
12'b10010011011100: data = 6'b111111;
12'b10010011011101: data = 6'b111111;
12'b10010011011110: data = 6'b111111;
12'b10010011011111: data = 6'b111111;
12'b10010011100000: data = 6'b111111;
12'b10010011100001: data = 6'b101010;
12'b10010011100010: data = 6'b101010;
12'b10010011100011: data = 6'b101010;
12'b10010011100100: data = 6'b101010;
12'b10010011100101: data = 6'b101010;
12'b10010011100110: data = 6'b101010;
12'b10010011100111: data = 6'b101010;
12'b10010011101000: data = 6'b101010;
12'b10010011101001: data = 6'b111111;
12'b10010011101010: data = 6'b111111;
12'b10010011101011: data = 6'b111111;
12'b10010011101100: data = 6'b111111;
12'b10010011101101: data = 6'b111111;
12'b10010011101110: data = 6'b111111;
12'b10010011101111: data = 6'b111111;
12'b10010011110000: data = 6'b111111;
12'b10010011110001: data = 6'b111111;
12'b10010011110010: data = 6'b111111;
12'b10010011110011: data = 6'b111111;
12'b10010011110100: data = 6'b111111;
12'b10010011110101: data = 6'b111111;
12'b10010011110110: data = 6'b111111;
12'b10010011110111: data = 6'b111111;
12'b10010011111000: data = 6'b111111;
12'b10010011111001: data = 6'b111111;
12'b10010011111010: data = 6'b111111;
12'b10010011111011: data = 6'b111111;
12'b10010011111100: data = 6'b111111;
12'b10010011111101: data = 6'b111111;
12'b10010011111110: data = 6'b111111;
12'b10010011111111: data = 6'b111111;
12'b100100110000000: data = 6'b111111;
12'b100100110000001: data = 6'b111111;
12'b100100110000010: data = 6'b111111;
12'b100100110000011: data = 6'b111111;
12'b100100110000100: data = 6'b101010;
12'b100100110000101: data = 6'b101010;
12'b100100110000110: data = 6'b101010;
12'b100100110000111: data = 6'b101010;
12'b100100110001000: data = 6'b101010;
12'b100100110001001: data = 6'b010101;
12'b100100110001010: data = 6'b010101;
12'b100100110001011: data = 6'b010101;
12'b100100110001100: data = 6'b000000;
12'b100100110001101: data = 6'b000000;
12'b100100110001110: data = 6'b101010;
12'b100100110001111: data = 6'b101010;
12'b100100110010000: data = 6'b101010;
12'b100100110010001: data = 6'b101010;
12'b100100110010010: data = 6'b010101;
12'b100100110010011: data = 6'b010101;
12'b100100110010100: data = 6'b010101;
12'b100100110010101: data = 6'b010101;
12'b100100110010110: data = 6'b010101;
12'b100100110010111: data = 6'b010101;
12'b100100110011000: data = 6'b010101;
12'b100100110011001: data = 6'b010101;
12'b100100110011010: data = 6'b010101;
12'b100100110011011: data = 6'b010101;
12'b100100110011100: data = 6'b010101;
12'b100100110011101: data = 6'b010101;
12'b100100110011110: data = 6'b010101;
12'b100100110011111: data = 6'b010101;
12'b100100110100000: data = 6'b010101;
12'b100100110100001: data = 6'b010101;
12'b100100110100010: data = 6'b010101;
12'b100100110100011: data = 6'b010101;
12'b100100110100100: data = 6'b010101;
12'b100100110100101: data = 6'b010101;
12'b100100110100110: data = 6'b010101;
12'b100100110100111: data = 6'b010101;
12'b100100110101000: data = 6'b010101;
12'b100100110101001: data = 6'b010101;
12'b100100110101010: data = 6'b010101;
12'b1001010000000: data = 6'b010101;
12'b1001010000001: data = 6'b010101;
12'b1001010000010: data = 6'b010101;
12'b1001010000011: data = 6'b010101;
12'b1001010000100: data = 6'b010101;
12'b1001010000101: data = 6'b010101;
12'b1001010000110: data = 6'b010101;
12'b1001010000111: data = 6'b010101;
12'b1001010001000: data = 6'b010101;
12'b1001010001001: data = 6'b010101;
12'b1001010001010: data = 6'b010101;
12'b1001010001011: data = 6'b010101;
12'b1001010001100: data = 6'b010101;
12'b1001010001101: data = 6'b010101;
12'b1001010001110: data = 6'b010101;
12'b1001010001111: data = 6'b010101;
12'b1001010010000: data = 6'b010101;
12'b1001010010001: data = 6'b010101;
12'b1001010010010: data = 6'b010101;
12'b1001010010011: data = 6'b010101;
12'b1001010010100: data = 6'b010101;
12'b1001010010101: data = 6'b010101;
12'b1001010010110: data = 6'b010101;
12'b1001010010111: data = 6'b010101;
12'b1001010011000: data = 6'b010101;
12'b1001010011001: data = 6'b101010;
12'b1001010011010: data = 6'b101010;
12'b1001010011011: data = 6'b101010;
12'b1001010011100: data = 6'b010101;
12'b1001010011101: data = 6'b000000;
12'b1001010011110: data = 6'b000000;
12'b1001010011111: data = 6'b010101;
12'b1001010100000: data = 6'b010101;
12'b1001010100001: data = 6'b010101;
12'b1001010100010: data = 6'b101010;
12'b1001010100011: data = 6'b101010;
12'b1001010100100: data = 6'b101010;
12'b1001010100101: data = 6'b101010;
12'b1001010100110: data = 6'b101010;
12'b1001010100111: data = 6'b111111;
12'b1001010101000: data = 6'b111111;
12'b1001010101001: data = 6'b111111;
12'b1001010101010: data = 6'b111111;
12'b1001010101011: data = 6'b111111;
12'b1001010101100: data = 6'b111111;
12'b1001010101101: data = 6'b111111;
12'b1001010101110: data = 6'b111111;
12'b1001010101111: data = 6'b111111;
12'b1001010110000: data = 6'b111111;
12'b1001010110001: data = 6'b111111;
12'b1001010110010: data = 6'b111111;
12'b1001010110011: data = 6'b111111;
12'b1001010110100: data = 6'b111111;
12'b1001010110101: data = 6'b111111;
12'b1001010110110: data = 6'b111111;
12'b1001010110111: data = 6'b111111;
12'b1001010111000: data = 6'b111111;
12'b1001010111001: data = 6'b111111;
12'b1001010111010: data = 6'b111111;
12'b1001010111011: data = 6'b111111;
12'b1001010111100: data = 6'b111111;
12'b1001010111101: data = 6'b111111;
12'b1001010111110: data = 6'b111111;
12'b1001010111111: data = 6'b111111;
12'b10010101000000: data = 6'b111111;
12'b10010101000001: data = 6'b111111;
12'b10010101000010: data = 6'b101010;
12'b10010101000011: data = 6'b101010;
12'b10010101000100: data = 6'b101010;
12'b10010101000101: data = 6'b101010;
12'b10010101000110: data = 6'b101010;
12'b10010101000111: data = 6'b101010;
12'b10010101001000: data = 6'b101010;
12'b10010101001001: data = 6'b101010;
12'b10010101001010: data = 6'b111111;
12'b10010101001011: data = 6'b111111;
12'b10010101001100: data = 6'b111111;
12'b10010101001101: data = 6'b111111;
12'b10010101001110: data = 6'b111111;
12'b10010101001111: data = 6'b111111;
12'b10010101010000: data = 6'b111111;
12'b10010101010001: data = 6'b111111;
12'b10010101010010: data = 6'b111111;
12'b10010101010011: data = 6'b111111;
12'b10010101010100: data = 6'b111111;
12'b10010101010101: data = 6'b111111;
12'b10010101010110: data = 6'b111111;
12'b10010101010111: data = 6'b111111;
12'b10010101011000: data = 6'b111111;
12'b10010101011001: data = 6'b111111;
12'b10010101011010: data = 6'b111111;
12'b10010101011011: data = 6'b111111;
12'b10010101011100: data = 6'b111111;
12'b10010101011101: data = 6'b111111;
12'b10010101011110: data = 6'b111111;
12'b10010101011111: data = 6'b111111;
12'b10010101100000: data = 6'b111111;
12'b10010101100001: data = 6'b101010;
12'b10010101100010: data = 6'b101001;
12'b10010101100011: data = 6'b101010;
12'b10010101100100: data = 6'b101010;
12'b10010101100101: data = 6'b101010;
12'b10010101100110: data = 6'b101010;
12'b10010101100111: data = 6'b101010;
12'b10010101101000: data = 6'b101010;
12'b10010101101001: data = 6'b111111;
12'b10010101101010: data = 6'b111111;
12'b10010101101011: data = 6'b111111;
12'b10010101101100: data = 6'b111111;
12'b10010101101101: data = 6'b111111;
12'b10010101101110: data = 6'b111111;
12'b10010101101111: data = 6'b111111;
12'b10010101110000: data = 6'b111111;
12'b10010101110001: data = 6'b111111;
12'b10010101110010: data = 6'b111111;
12'b10010101110011: data = 6'b111111;
12'b10010101110100: data = 6'b111111;
12'b10010101110101: data = 6'b111111;
12'b10010101110110: data = 6'b111111;
12'b10010101110111: data = 6'b111111;
12'b10010101111000: data = 6'b111111;
12'b10010101111001: data = 6'b111111;
12'b10010101111010: data = 6'b111111;
12'b10010101111011: data = 6'b111111;
12'b10010101111100: data = 6'b111111;
12'b10010101111101: data = 6'b111111;
12'b10010101111110: data = 6'b111111;
12'b10010101111111: data = 6'b111111;
12'b100101010000000: data = 6'b111111;
12'b100101010000001: data = 6'b111111;
12'b100101010000010: data = 6'b111111;
12'b100101010000011: data = 6'b111111;
12'b100101010000100: data = 6'b101010;
12'b100101010000101: data = 6'b101010;
12'b100101010000110: data = 6'b101010;
12'b100101010000111: data = 6'b101010;
12'b100101010001000: data = 6'b101010;
12'b100101010001001: data = 6'b010101;
12'b100101010001010: data = 6'b010101;
12'b100101010001011: data = 6'b010101;
12'b100101010001100: data = 6'b000000;
12'b100101010001101: data = 6'b000000;
12'b100101010001110: data = 6'b101010;
12'b100101010001111: data = 6'b101010;
12'b100101010010000: data = 6'b101010;
12'b100101010010001: data = 6'b101010;
12'b100101010010010: data = 6'b010101;
12'b100101010010011: data = 6'b010101;
12'b100101010010100: data = 6'b010101;
12'b100101010010101: data = 6'b010101;
12'b100101010010110: data = 6'b010101;
12'b100101010010111: data = 6'b010101;
12'b100101010011000: data = 6'b010101;
12'b100101010011001: data = 6'b010101;
12'b100101010011010: data = 6'b010101;
12'b100101010011011: data = 6'b010101;
12'b100101010011100: data = 6'b010101;
12'b100101010011101: data = 6'b010101;
12'b100101010011110: data = 6'b010101;
12'b100101010011111: data = 6'b010101;
12'b100101010100000: data = 6'b010101;
12'b100101010100001: data = 6'b010101;
12'b100101010100010: data = 6'b010101;
12'b100101010100011: data = 6'b010101;
12'b100101010100100: data = 6'b010101;
12'b100101010100101: data = 6'b010101;
12'b100101010100110: data = 6'b010101;
12'b100101010100111: data = 6'b010101;
12'b100101010101000: data = 6'b010101;
12'b100101010101001: data = 6'b010101;
12'b100101010101010: data = 6'b010101;
12'b1001011000000: data = 6'b010101;
12'b1001011000001: data = 6'b010101;
12'b1001011000010: data = 6'b010101;
12'b1001011000011: data = 6'b010101;
12'b1001011000100: data = 6'b010101;
12'b1001011000101: data = 6'b010101;
12'b1001011000110: data = 6'b010101;
12'b1001011000111: data = 6'b010101;
12'b1001011001000: data = 6'b010101;
12'b1001011001001: data = 6'b010101;
12'b1001011001010: data = 6'b010101;
12'b1001011001011: data = 6'b010101;
12'b1001011001100: data = 6'b010101;
12'b1001011001101: data = 6'b010101;
12'b1001011001110: data = 6'b010101;
12'b1001011001111: data = 6'b010101;
12'b1001011010000: data = 6'b010101;
12'b1001011010001: data = 6'b010101;
12'b1001011010010: data = 6'b010101;
12'b1001011010011: data = 6'b010101;
12'b1001011010100: data = 6'b010101;
12'b1001011010101: data = 6'b010101;
12'b1001011010110: data = 6'b010101;
12'b1001011010111: data = 6'b010101;
12'b1001011011000: data = 6'b010101;
12'b1001011011001: data = 6'b101010;
12'b1001011011010: data = 6'b101010;
12'b1001011011011: data = 6'b101010;
12'b1001011011100: data = 6'b010101;
12'b1001011011101: data = 6'b000000;
12'b1001011011110: data = 6'b000000;
12'b1001011011111: data = 6'b010101;
12'b1001011100000: data = 6'b010101;
12'b1001011100001: data = 6'b010101;
12'b1001011100010: data = 6'b101010;
12'b1001011100011: data = 6'b101010;
12'b1001011100100: data = 6'b101010;
12'b1001011100101: data = 6'b101010;
12'b1001011100110: data = 6'b101010;
12'b1001011100111: data = 6'b111111;
12'b1001011101000: data = 6'b111111;
12'b1001011101001: data = 6'b111111;
12'b1001011101010: data = 6'b111111;
12'b1001011101011: data = 6'b111111;
12'b1001011101100: data = 6'b111111;
12'b1001011101101: data = 6'b111111;
12'b1001011101110: data = 6'b111111;
12'b1001011101111: data = 6'b111111;
12'b1001011110000: data = 6'b111111;
12'b1001011110001: data = 6'b111111;
12'b1001011110010: data = 6'b111111;
12'b1001011110011: data = 6'b111111;
12'b1001011110100: data = 6'b111111;
12'b1001011110101: data = 6'b111111;
12'b1001011110110: data = 6'b111111;
12'b1001011110111: data = 6'b111111;
12'b1001011111000: data = 6'b111111;
12'b1001011111001: data = 6'b111111;
12'b1001011111010: data = 6'b111111;
12'b1001011111011: data = 6'b111111;
12'b1001011111100: data = 6'b111111;
12'b1001011111101: data = 6'b111111;
12'b1001011111110: data = 6'b111111;
12'b1001011111111: data = 6'b111111;
12'b10010111000000: data = 6'b111111;
12'b10010111000001: data = 6'b111111;
12'b10010111000010: data = 6'b101010;
12'b10010111000011: data = 6'b101010;
12'b10010111000100: data = 6'b101010;
12'b10010111000101: data = 6'b101010;
12'b10010111000110: data = 6'b101010;
12'b10010111000111: data = 6'b101010;
12'b10010111001000: data = 6'b101001;
12'b10010111001001: data = 6'b101010;
12'b10010111001010: data = 6'b111111;
12'b10010111001011: data = 6'b111111;
12'b10010111001100: data = 6'b111111;
12'b10010111001101: data = 6'b111111;
12'b10010111001110: data = 6'b111111;
12'b10010111001111: data = 6'b111111;
12'b10010111010000: data = 6'b111111;
12'b10010111010001: data = 6'b111111;
12'b10010111010010: data = 6'b111111;
12'b10010111010011: data = 6'b111111;
12'b10010111010100: data = 6'b111111;
12'b10010111010101: data = 6'b111111;
12'b10010111010110: data = 6'b111111;
12'b10010111010111: data = 6'b111111;
12'b10010111011000: data = 6'b111111;
12'b10010111011001: data = 6'b111111;
12'b10010111011010: data = 6'b111111;
12'b10010111011011: data = 6'b111111;
12'b10010111011100: data = 6'b111111;
12'b10010111011101: data = 6'b111111;
12'b10010111011110: data = 6'b111111;
12'b10010111011111: data = 6'b111111;
12'b10010111100000: data = 6'b111111;
12'b10010111100001: data = 6'b101010;
12'b10010111100010: data = 6'b010101;
12'b10010111100011: data = 6'b101001;
12'b10010111100100: data = 6'b101010;
12'b10010111100101: data = 6'b101010;
12'b10010111100110: data = 6'b101010;
12'b10010111100111: data = 6'b101010;
12'b10010111101000: data = 6'b101010;
12'b10010111101001: data = 6'b111111;
12'b10010111101010: data = 6'b111111;
12'b10010111101011: data = 6'b111111;
12'b10010111101100: data = 6'b111111;
12'b10010111101101: data = 6'b111111;
12'b10010111101110: data = 6'b111111;
12'b10010111101111: data = 6'b111111;
12'b10010111110000: data = 6'b111111;
12'b10010111110001: data = 6'b111111;
12'b10010111110010: data = 6'b111111;
12'b10010111110011: data = 6'b111111;
12'b10010111110100: data = 6'b111111;
12'b10010111110101: data = 6'b111111;
12'b10010111110110: data = 6'b111111;
12'b10010111110111: data = 6'b111111;
12'b10010111111000: data = 6'b111111;
12'b10010111111001: data = 6'b111111;
12'b10010111111010: data = 6'b111111;
12'b10010111111011: data = 6'b111111;
12'b10010111111100: data = 6'b111111;
12'b10010111111101: data = 6'b111111;
12'b10010111111110: data = 6'b111111;
12'b10010111111111: data = 6'b111111;
12'b100101110000000: data = 6'b111111;
12'b100101110000001: data = 6'b111111;
12'b100101110000010: data = 6'b111111;
12'b100101110000011: data = 6'b111111;
12'b100101110000100: data = 6'b101010;
12'b100101110000101: data = 6'b101010;
12'b100101110000110: data = 6'b101010;
12'b100101110000111: data = 6'b101010;
12'b100101110001000: data = 6'b101010;
12'b100101110001001: data = 6'b010101;
12'b100101110001010: data = 6'b010101;
12'b100101110001011: data = 6'b010101;
12'b100101110001100: data = 6'b000000;
12'b100101110001101: data = 6'b000000;
12'b100101110001110: data = 6'b101010;
12'b100101110001111: data = 6'b101010;
12'b100101110010000: data = 6'b101010;
12'b100101110010001: data = 6'b101010;
12'b100101110010010: data = 6'b010101;
12'b100101110010011: data = 6'b010101;
12'b100101110010100: data = 6'b010101;
12'b100101110010101: data = 6'b010101;
12'b100101110010110: data = 6'b010101;
12'b100101110010111: data = 6'b010101;
12'b100101110011000: data = 6'b010101;
12'b100101110011001: data = 6'b010101;
12'b100101110011010: data = 6'b010101;
12'b100101110011011: data = 6'b010101;
12'b100101110011100: data = 6'b010101;
12'b100101110011101: data = 6'b010101;
12'b100101110011110: data = 6'b010101;
12'b100101110011111: data = 6'b010101;
12'b100101110100000: data = 6'b010101;
12'b100101110100001: data = 6'b010101;
12'b100101110100010: data = 6'b010101;
12'b100101110100011: data = 6'b010101;
12'b100101110100100: data = 6'b010101;
12'b100101110100101: data = 6'b010101;
12'b100101110100110: data = 6'b010101;
12'b100101110100111: data = 6'b010101;
12'b100101110101000: data = 6'b010101;
12'b100101110101001: data = 6'b010101;
12'b100101110101010: data = 6'b010101;
12'b1001100000000: data = 6'b010101;
12'b1001100000001: data = 6'b010101;
12'b1001100000010: data = 6'b010101;
12'b1001100000011: data = 6'b010101;
12'b1001100000100: data = 6'b010101;
12'b1001100000101: data = 6'b010101;
12'b1001100000110: data = 6'b010101;
12'b1001100000111: data = 6'b010101;
12'b1001100001000: data = 6'b010101;
12'b1001100001001: data = 6'b010101;
12'b1001100001010: data = 6'b010101;
12'b1001100001011: data = 6'b010101;
12'b1001100001100: data = 6'b010101;
12'b1001100001101: data = 6'b010101;
12'b1001100001110: data = 6'b010101;
12'b1001100001111: data = 6'b010101;
12'b1001100010000: data = 6'b010101;
12'b1001100010001: data = 6'b010101;
12'b1001100010010: data = 6'b010101;
12'b1001100010011: data = 6'b010101;
12'b1001100010100: data = 6'b010101;
12'b1001100010101: data = 6'b010101;
12'b1001100010110: data = 6'b010101;
12'b1001100010111: data = 6'b010101;
12'b1001100011000: data = 6'b010101;
12'b1001100011001: data = 6'b101010;
12'b1001100011010: data = 6'b101010;
12'b1001100011011: data = 6'b101010;
12'b1001100011100: data = 6'b010101;
12'b1001100011101: data = 6'b000000;
12'b1001100011110: data = 6'b000000;
12'b1001100011111: data = 6'b010101;
12'b1001100100000: data = 6'b010101;
12'b1001100100001: data = 6'b010101;
12'b1001100100010: data = 6'b101010;
12'b1001100100011: data = 6'b101010;
12'b1001100100100: data = 6'b101010;
12'b1001100100101: data = 6'b101010;
12'b1001100100110: data = 6'b101010;
12'b1001100100111: data = 6'b111111;
12'b1001100101000: data = 6'b111111;
12'b1001100101001: data = 6'b111111;
12'b1001100101010: data = 6'b111111;
12'b1001100101011: data = 6'b111111;
12'b1001100101100: data = 6'b111111;
12'b1001100101101: data = 6'b111111;
12'b1001100101110: data = 6'b111111;
12'b1001100101111: data = 6'b111111;
12'b1001100110000: data = 6'b111111;
12'b1001100110001: data = 6'b111111;
12'b1001100110010: data = 6'b111111;
12'b1001100110011: data = 6'b111111;
12'b1001100110100: data = 6'b111111;
12'b1001100110101: data = 6'b111111;
12'b1001100110110: data = 6'b111111;
12'b1001100110111: data = 6'b111111;
12'b1001100111000: data = 6'b111111;
12'b1001100111001: data = 6'b111111;
12'b1001100111010: data = 6'b111111;
12'b1001100111011: data = 6'b111111;
12'b1001100111100: data = 6'b111111;
12'b1001100111101: data = 6'b111111;
12'b1001100111110: data = 6'b111111;
12'b1001100111111: data = 6'b111111;
12'b10011001000000: data = 6'b111111;
12'b10011001000001: data = 6'b111111;
12'b10011001000010: data = 6'b101010;
12'b10011001000011: data = 6'b101010;
12'b10011001000100: data = 6'b101010;
12'b10011001000101: data = 6'b101010;
12'b10011001000110: data = 6'b101010;
12'b10011001000111: data = 6'b101010;
12'b10011001001000: data = 6'b010101;
12'b10011001001001: data = 6'b101010;
12'b10011001001010: data = 6'b111111;
12'b10011001001011: data = 6'b111111;
12'b10011001001100: data = 6'b111111;
12'b10011001001101: data = 6'b111111;
12'b10011001001110: data = 6'b111111;
12'b10011001001111: data = 6'b111111;
12'b10011001010000: data = 6'b111111;
12'b10011001010001: data = 6'b111111;
12'b10011001010010: data = 6'b111111;
12'b10011001010011: data = 6'b111111;
12'b10011001010100: data = 6'b111111;
12'b10011001010101: data = 6'b111111;
12'b10011001010110: data = 6'b111111;
12'b10011001010111: data = 6'b111111;
12'b10011001011000: data = 6'b111111;
12'b10011001011001: data = 6'b111111;
12'b10011001011010: data = 6'b111111;
12'b10011001011011: data = 6'b111111;
12'b10011001011100: data = 6'b111111;
12'b10011001011101: data = 6'b111111;
12'b10011001011110: data = 6'b111111;
12'b10011001011111: data = 6'b111111;
12'b10011001100000: data = 6'b111111;
12'b10011001100001: data = 6'b101010;
12'b10011001100010: data = 6'b010101;
12'b10011001100011: data = 6'b101001;
12'b10011001100100: data = 6'b101010;
12'b10011001100101: data = 6'b101010;
12'b10011001100110: data = 6'b101010;
12'b10011001100111: data = 6'b101010;
12'b10011001101000: data = 6'b101010;
12'b10011001101001: data = 6'b111111;
12'b10011001101010: data = 6'b111111;
12'b10011001101011: data = 6'b111111;
12'b10011001101100: data = 6'b111111;
12'b10011001101101: data = 6'b111111;
12'b10011001101110: data = 6'b111111;
12'b10011001101111: data = 6'b111111;
12'b10011001110000: data = 6'b111111;
12'b10011001110001: data = 6'b111111;
12'b10011001110010: data = 6'b111111;
12'b10011001110011: data = 6'b111111;
12'b10011001110100: data = 6'b111111;
12'b10011001110101: data = 6'b111111;
12'b10011001110110: data = 6'b111111;
12'b10011001110111: data = 6'b111111;
12'b10011001111000: data = 6'b111111;
12'b10011001111001: data = 6'b111111;
12'b10011001111010: data = 6'b111111;
12'b10011001111011: data = 6'b111111;
12'b10011001111100: data = 6'b111111;
12'b10011001111101: data = 6'b111111;
12'b10011001111110: data = 6'b111111;
12'b10011001111111: data = 6'b111111;
12'b100110010000000: data = 6'b111111;
12'b100110010000001: data = 6'b111111;
12'b100110010000010: data = 6'b111111;
12'b100110010000011: data = 6'b111111;
12'b100110010000100: data = 6'b101010;
12'b100110010000101: data = 6'b101010;
12'b100110010000110: data = 6'b101010;
12'b100110010000111: data = 6'b101010;
12'b100110010001000: data = 6'b101010;
12'b100110010001001: data = 6'b010101;
12'b100110010001010: data = 6'b010101;
12'b100110010001011: data = 6'b010101;
12'b100110010001100: data = 6'b000000;
12'b100110010001101: data = 6'b000000;
12'b100110010001110: data = 6'b101010;
12'b100110010001111: data = 6'b101010;
12'b100110010010000: data = 6'b101010;
12'b100110010010001: data = 6'b101010;
12'b100110010010010: data = 6'b010101;
12'b100110010010011: data = 6'b010101;
12'b100110010010100: data = 6'b010101;
12'b100110010010101: data = 6'b010101;
12'b100110010010110: data = 6'b010101;
12'b100110010010111: data = 6'b010101;
12'b100110010011000: data = 6'b010101;
12'b100110010011001: data = 6'b010101;
12'b100110010011010: data = 6'b010101;
12'b100110010011011: data = 6'b010101;
12'b100110010011100: data = 6'b010101;
12'b100110010011101: data = 6'b010101;
12'b100110010011110: data = 6'b010101;
12'b100110010011111: data = 6'b010101;
12'b100110010100000: data = 6'b010101;
12'b100110010100001: data = 6'b010101;
12'b100110010100010: data = 6'b010101;
12'b100110010100011: data = 6'b010101;
12'b100110010100100: data = 6'b010101;
12'b100110010100101: data = 6'b010101;
12'b100110010100110: data = 6'b010101;
12'b100110010100111: data = 6'b010101;
12'b100110010101000: data = 6'b010101;
12'b100110010101001: data = 6'b010101;
12'b100110010101010: data = 6'b010101;
12'b1001101000000: data = 6'b010101;
12'b1001101000001: data = 6'b010101;
12'b1001101000010: data = 6'b010101;
12'b1001101000011: data = 6'b010101;
12'b1001101000100: data = 6'b010101;
12'b1001101000101: data = 6'b010101;
12'b1001101000110: data = 6'b010101;
12'b1001101000111: data = 6'b010101;
12'b1001101001000: data = 6'b010101;
12'b1001101001001: data = 6'b010101;
12'b1001101001010: data = 6'b010101;
12'b1001101001011: data = 6'b010101;
12'b1001101001100: data = 6'b010101;
12'b1001101001101: data = 6'b010101;
12'b1001101001110: data = 6'b010101;
12'b1001101001111: data = 6'b010101;
12'b1001101010000: data = 6'b010101;
12'b1001101010001: data = 6'b010101;
12'b1001101010010: data = 6'b010101;
12'b1001101010011: data = 6'b010101;
12'b1001101010100: data = 6'b010101;
12'b1001101010101: data = 6'b010101;
12'b1001101010110: data = 6'b010101;
12'b1001101010111: data = 6'b010101;
12'b1001101011000: data = 6'b010101;
12'b1001101011001: data = 6'b101010;
12'b1001101011010: data = 6'b101010;
12'b1001101011011: data = 6'b101010;
12'b1001101011100: data = 6'b010101;
12'b1001101011101: data = 6'b000000;
12'b1001101011110: data = 6'b000000;
12'b1001101011111: data = 6'b010101;
12'b1001101100000: data = 6'b010101;
12'b1001101100001: data = 6'b010101;
12'b1001101100010: data = 6'b101010;
12'b1001101100011: data = 6'b101010;
12'b1001101100100: data = 6'b101010;
12'b1001101100101: data = 6'b101010;
12'b1001101100110: data = 6'b101010;
12'b1001101100111: data = 6'b111111;
12'b1001101101000: data = 6'b111111;
12'b1001101101001: data = 6'b111111;
12'b1001101101010: data = 6'b111111;
12'b1001101101011: data = 6'b111111;
12'b1001101101100: data = 6'b111111;
12'b1001101101101: data = 6'b111111;
12'b1001101101110: data = 6'b111111;
12'b1001101101111: data = 6'b111111;
12'b1001101110000: data = 6'b111111;
12'b1001101110001: data = 6'b111111;
12'b1001101110010: data = 6'b111111;
12'b1001101110011: data = 6'b111111;
12'b1001101110100: data = 6'b111111;
12'b1001101110101: data = 6'b111111;
12'b1001101110110: data = 6'b111111;
12'b1001101110111: data = 6'b111111;
12'b1001101111000: data = 6'b111111;
12'b1001101111001: data = 6'b111111;
12'b1001101111010: data = 6'b111111;
12'b1001101111011: data = 6'b111111;
12'b1001101111100: data = 6'b111111;
12'b1001101111101: data = 6'b111111;
12'b1001101111110: data = 6'b111111;
12'b1001101111111: data = 6'b111111;
12'b10011011000000: data = 6'b111111;
12'b10011011000001: data = 6'b111111;
12'b10011011000010: data = 6'b101010;
12'b10011011000011: data = 6'b101010;
12'b10011011000100: data = 6'b101010;
12'b10011011000101: data = 6'b101010;
12'b10011011000110: data = 6'b101010;
12'b10011011000111: data = 6'b101010;
12'b10011011001000: data = 6'b010101;
12'b10011011001001: data = 6'b101010;
12'b10011011001010: data = 6'b111111;
12'b10011011001011: data = 6'b111111;
12'b10011011001100: data = 6'b111111;
12'b10011011001101: data = 6'b111111;
12'b10011011001110: data = 6'b111111;
12'b10011011001111: data = 6'b111111;
12'b10011011010000: data = 6'b111111;
12'b10011011010001: data = 6'b111111;
12'b10011011010010: data = 6'b111111;
12'b10011011010011: data = 6'b111111;
12'b10011011010100: data = 6'b111111;
12'b10011011010101: data = 6'b111111;
12'b10011011010110: data = 6'b111111;
12'b10011011010111: data = 6'b111111;
12'b10011011011000: data = 6'b111111;
12'b10011011011001: data = 6'b111111;
12'b10011011011010: data = 6'b111111;
12'b10011011011011: data = 6'b111111;
12'b10011011011100: data = 6'b111111;
12'b10011011011101: data = 6'b111111;
12'b10011011011110: data = 6'b111111;
12'b10011011011111: data = 6'b111111;
12'b10011011100000: data = 6'b111111;
12'b10011011100001: data = 6'b101010;
12'b10011011100010: data = 6'b010101;
12'b10011011100011: data = 6'b101001;
12'b10011011100100: data = 6'b101010;
12'b10011011100101: data = 6'b101010;
12'b10011011100110: data = 6'b101010;
12'b10011011100111: data = 6'b101010;
12'b10011011101000: data = 6'b101010;
12'b10011011101001: data = 6'b111111;
12'b10011011101010: data = 6'b111111;
12'b10011011101011: data = 6'b111111;
12'b10011011101100: data = 6'b111111;
12'b10011011101101: data = 6'b111111;
12'b10011011101110: data = 6'b111111;
12'b10011011101111: data = 6'b111111;
12'b10011011110000: data = 6'b111111;
12'b10011011110001: data = 6'b111111;
12'b10011011110010: data = 6'b111111;
12'b10011011110011: data = 6'b111111;
12'b10011011110100: data = 6'b111111;
12'b10011011110101: data = 6'b111111;
12'b10011011110110: data = 6'b111111;
12'b10011011110111: data = 6'b111111;
12'b10011011111000: data = 6'b111111;
12'b10011011111001: data = 6'b111111;
12'b10011011111010: data = 6'b111111;
12'b10011011111011: data = 6'b111111;
12'b10011011111100: data = 6'b111111;
12'b10011011111101: data = 6'b111111;
12'b10011011111110: data = 6'b111111;
12'b10011011111111: data = 6'b111111;
12'b100110110000000: data = 6'b111111;
12'b100110110000001: data = 6'b111111;
12'b100110110000010: data = 6'b111111;
12'b100110110000011: data = 6'b111111;
12'b100110110000100: data = 6'b101010;
12'b100110110000101: data = 6'b101010;
12'b100110110000110: data = 6'b101010;
12'b100110110000111: data = 6'b101010;
12'b100110110001000: data = 6'b101010;
12'b100110110001001: data = 6'b010101;
12'b100110110001010: data = 6'b010101;
12'b100110110001011: data = 6'b010101;
12'b100110110001100: data = 6'b000000;
12'b100110110001101: data = 6'b000000;
12'b100110110001110: data = 6'b101010;
12'b100110110001111: data = 6'b101010;
12'b100110110010000: data = 6'b101010;
12'b100110110010001: data = 6'b101010;
12'b100110110010010: data = 6'b010101;
12'b100110110010011: data = 6'b010101;
12'b100110110010100: data = 6'b010101;
12'b100110110010101: data = 6'b010101;
12'b100110110010110: data = 6'b010101;
12'b100110110010111: data = 6'b010101;
12'b100110110011000: data = 6'b010101;
12'b100110110011001: data = 6'b010101;
12'b100110110011010: data = 6'b010101;
12'b100110110011011: data = 6'b010101;
12'b100110110011100: data = 6'b010101;
12'b100110110011101: data = 6'b010101;
12'b100110110011110: data = 6'b010101;
12'b100110110011111: data = 6'b010101;
12'b100110110100000: data = 6'b010101;
12'b100110110100001: data = 6'b010101;
12'b100110110100010: data = 6'b010101;
12'b100110110100011: data = 6'b010101;
12'b100110110100100: data = 6'b010101;
12'b100110110100101: data = 6'b010101;
12'b100110110100110: data = 6'b010101;
12'b100110110100111: data = 6'b010101;
12'b100110110101000: data = 6'b010101;
12'b100110110101001: data = 6'b010101;
12'b100110110101010: data = 6'b010101;
12'b1001110000000: data = 6'b010101;
12'b1001110000001: data = 6'b010101;
12'b1001110000010: data = 6'b010101;
12'b1001110000011: data = 6'b010101;
12'b1001110000100: data = 6'b010101;
12'b1001110000101: data = 6'b010101;
12'b1001110000110: data = 6'b010101;
12'b1001110000111: data = 6'b010101;
12'b1001110001000: data = 6'b010101;
12'b1001110001001: data = 6'b010101;
12'b1001110001010: data = 6'b010101;
12'b1001110001011: data = 6'b010101;
12'b1001110001100: data = 6'b010101;
12'b1001110001101: data = 6'b010101;
12'b1001110001110: data = 6'b010101;
12'b1001110001111: data = 6'b010101;
12'b1001110010000: data = 6'b010101;
12'b1001110010001: data = 6'b010101;
12'b1001110010010: data = 6'b010101;
12'b1001110010011: data = 6'b010101;
12'b1001110010100: data = 6'b010101;
12'b1001110010101: data = 6'b010101;
12'b1001110010110: data = 6'b010101;
12'b1001110010111: data = 6'b010101;
12'b1001110011000: data = 6'b010101;
12'b1001110011001: data = 6'b101010;
12'b1001110011010: data = 6'b101010;
12'b1001110011011: data = 6'b101010;
12'b1001110011100: data = 6'b010101;
12'b1001110011101: data = 6'b000000;
12'b1001110011110: data = 6'b000000;
12'b1001110011111: data = 6'b010101;
12'b1001110100000: data = 6'b010101;
12'b1001110100001: data = 6'b010101;
12'b1001110100010: data = 6'b101010;
12'b1001110100011: data = 6'b101010;
12'b1001110100100: data = 6'b101010;
12'b1001110100101: data = 6'b101010;
12'b1001110100110: data = 6'b101010;
12'b1001110100111: data = 6'b111111;
12'b1001110101000: data = 6'b111111;
12'b1001110101001: data = 6'b111111;
12'b1001110101010: data = 6'b111111;
12'b1001110101011: data = 6'b111111;
12'b1001110101100: data = 6'b111111;
12'b1001110101101: data = 6'b111111;
12'b1001110101110: data = 6'b111111;
12'b1001110101111: data = 6'b111111;
12'b1001110110000: data = 6'b111111;
12'b1001110110001: data = 6'b111111;
12'b1001110110010: data = 6'b111111;
12'b1001110110011: data = 6'b111111;
12'b1001110110100: data = 6'b111111;
12'b1001110110101: data = 6'b111111;
12'b1001110110110: data = 6'b111111;
12'b1001110110111: data = 6'b111111;
12'b1001110111000: data = 6'b111111;
12'b1001110111001: data = 6'b111111;
12'b1001110111010: data = 6'b111111;
12'b1001110111011: data = 6'b111111;
12'b1001110111100: data = 6'b111111;
12'b1001110111101: data = 6'b111111;
12'b1001110111110: data = 6'b111111;
12'b1001110111111: data = 6'b111111;
12'b10011101000000: data = 6'b111111;
12'b10011101000001: data = 6'b111111;
12'b10011101000010: data = 6'b101010;
12'b10011101000011: data = 6'b101010;
12'b10011101000100: data = 6'b101010;
12'b10011101000101: data = 6'b101010;
12'b10011101000110: data = 6'b101010;
12'b10011101000111: data = 6'b101010;
12'b10011101001000: data = 6'b010101;
12'b10011101001001: data = 6'b101010;
12'b10011101001010: data = 6'b111111;
12'b10011101001011: data = 6'b111111;
12'b10011101001100: data = 6'b111111;
12'b10011101001101: data = 6'b111111;
12'b10011101001110: data = 6'b111111;
12'b10011101001111: data = 6'b111111;
12'b10011101010000: data = 6'b111111;
12'b10011101010001: data = 6'b111111;
12'b10011101010010: data = 6'b111111;
12'b10011101010011: data = 6'b111111;
12'b10011101010100: data = 6'b111111;
12'b10011101010101: data = 6'b111111;
12'b10011101010110: data = 6'b111111;
12'b10011101010111: data = 6'b111111;
12'b10011101011000: data = 6'b111111;
12'b10011101011001: data = 6'b111111;
12'b10011101011010: data = 6'b111111;
12'b10011101011011: data = 6'b111111;
12'b10011101011100: data = 6'b111111;
12'b10011101011101: data = 6'b111111;
12'b10011101011110: data = 6'b111111;
12'b10011101011111: data = 6'b111111;
12'b10011101100000: data = 6'b111111;
12'b10011101100001: data = 6'b101010;
12'b10011101100010: data = 6'b010101;
12'b10011101100011: data = 6'b101001;
12'b10011101100100: data = 6'b101010;
12'b10011101100101: data = 6'b101010;
12'b10011101100110: data = 6'b101010;
12'b10011101100111: data = 6'b101010;
12'b10011101101000: data = 6'b101010;
12'b10011101101001: data = 6'b111111;
12'b10011101101010: data = 6'b111111;
12'b10011101101011: data = 6'b111111;
12'b10011101101100: data = 6'b111111;
12'b10011101101101: data = 6'b111111;
12'b10011101101110: data = 6'b111111;
12'b10011101101111: data = 6'b111111;
12'b10011101110000: data = 6'b111111;
12'b10011101110001: data = 6'b111111;
12'b10011101110010: data = 6'b111111;
12'b10011101110011: data = 6'b111111;
12'b10011101110100: data = 6'b111111;
12'b10011101110101: data = 6'b111111;
12'b10011101110110: data = 6'b111111;
12'b10011101110111: data = 6'b111111;
12'b10011101111000: data = 6'b111111;
12'b10011101111001: data = 6'b111111;
12'b10011101111010: data = 6'b111111;
12'b10011101111011: data = 6'b111111;
12'b10011101111100: data = 6'b111111;
12'b10011101111101: data = 6'b111111;
12'b10011101111110: data = 6'b111111;
12'b10011101111111: data = 6'b111111;
12'b100111010000000: data = 6'b111111;
12'b100111010000001: data = 6'b111111;
12'b100111010000010: data = 6'b111111;
12'b100111010000011: data = 6'b111111;
12'b100111010000100: data = 6'b101010;
12'b100111010000101: data = 6'b101010;
12'b100111010000110: data = 6'b101010;
12'b100111010000111: data = 6'b101010;
12'b100111010001000: data = 6'b101010;
12'b100111010001001: data = 6'b010101;
12'b100111010001010: data = 6'b010101;
12'b100111010001011: data = 6'b010101;
12'b100111010001100: data = 6'b000000;
12'b100111010001101: data = 6'b000000;
12'b100111010001110: data = 6'b101010;
12'b100111010001111: data = 6'b101010;
12'b100111010010000: data = 6'b101010;
12'b100111010010001: data = 6'b101010;
12'b100111010010010: data = 6'b010101;
12'b100111010010011: data = 6'b010101;
12'b100111010010100: data = 6'b010101;
12'b100111010010101: data = 6'b010101;
12'b100111010010110: data = 6'b010101;
12'b100111010010111: data = 6'b010101;
12'b100111010011000: data = 6'b010101;
12'b100111010011001: data = 6'b010101;
12'b100111010011010: data = 6'b010101;
12'b100111010011011: data = 6'b010101;
12'b100111010011100: data = 6'b010101;
12'b100111010011101: data = 6'b010101;
12'b100111010011110: data = 6'b010101;
12'b100111010011111: data = 6'b010101;
12'b100111010100000: data = 6'b010101;
12'b100111010100001: data = 6'b010101;
12'b100111010100010: data = 6'b010101;
12'b100111010100011: data = 6'b010101;
12'b100111010100100: data = 6'b010101;
12'b100111010100101: data = 6'b010101;
12'b100111010100110: data = 6'b010101;
12'b100111010100111: data = 6'b010101;
12'b100111010101000: data = 6'b010101;
12'b100111010101001: data = 6'b010101;
12'b100111010101010: data = 6'b010101;
12'b1001111000000: data = 6'b010101;
12'b1001111000001: data = 6'b010101;
12'b1001111000010: data = 6'b010101;
12'b1001111000011: data = 6'b010101;
12'b1001111000100: data = 6'b010101;
12'b1001111000101: data = 6'b010101;
12'b1001111000110: data = 6'b010101;
12'b1001111000111: data = 6'b010101;
12'b1001111001000: data = 6'b010101;
12'b1001111001001: data = 6'b010101;
12'b1001111001010: data = 6'b010101;
12'b1001111001011: data = 6'b010101;
12'b1001111001100: data = 6'b010101;
12'b1001111001101: data = 6'b010101;
12'b1001111001110: data = 6'b010101;
12'b1001111001111: data = 6'b010101;
12'b1001111010000: data = 6'b010101;
12'b1001111010001: data = 6'b010101;
12'b1001111010010: data = 6'b010101;
12'b1001111010011: data = 6'b010101;
12'b1001111010100: data = 6'b010101;
12'b1001111010101: data = 6'b010101;
12'b1001111010110: data = 6'b010101;
12'b1001111010111: data = 6'b010101;
12'b1001111011000: data = 6'b010101;
12'b1001111011001: data = 6'b101010;
12'b1001111011010: data = 6'b101010;
12'b1001111011011: data = 6'b101010;
12'b1001111011100: data = 6'b010101;
12'b1001111011101: data = 6'b000000;
12'b1001111011110: data = 6'b000000;
12'b1001111011111: data = 6'b010101;
12'b1001111100000: data = 6'b010101;
12'b1001111100001: data = 6'b010101;
12'b1001111100010: data = 6'b101010;
12'b1001111100011: data = 6'b101010;
12'b1001111100100: data = 6'b101010;
12'b1001111100101: data = 6'b101010;
12'b1001111100110: data = 6'b101010;
12'b1001111100111: data = 6'b111111;
12'b1001111101000: data = 6'b111111;
12'b1001111101001: data = 6'b111111;
12'b1001111101010: data = 6'b111111;
12'b1001111101011: data = 6'b111111;
12'b1001111101100: data = 6'b111111;
12'b1001111101101: data = 6'b111111;
12'b1001111101110: data = 6'b111111;
12'b1001111101111: data = 6'b111111;
12'b1001111110000: data = 6'b111111;
12'b1001111110001: data = 6'b111111;
12'b1001111110010: data = 6'b111111;
12'b1001111110011: data = 6'b111111;
12'b1001111110100: data = 6'b111111;
12'b1001111110101: data = 6'b111111;
12'b1001111110110: data = 6'b111111;
12'b1001111110111: data = 6'b111111;
12'b1001111111000: data = 6'b111111;
12'b1001111111001: data = 6'b111111;
12'b1001111111010: data = 6'b111111;
12'b1001111111011: data = 6'b111111;
12'b1001111111100: data = 6'b111111;
12'b1001111111101: data = 6'b111111;
12'b1001111111110: data = 6'b111111;
12'b1001111111111: data = 6'b111111;
12'b10011111000000: data = 6'b111111;
12'b10011111000001: data = 6'b111111;
12'b10011111000010: data = 6'b101010;
12'b10011111000011: data = 6'b101010;
12'b10011111000100: data = 6'b101010;
12'b10011111000101: data = 6'b101010;
12'b10011111000110: data = 6'b101010;
12'b10011111000111: data = 6'b101010;
12'b10011111001000: data = 6'b010101;
12'b10011111001001: data = 6'b101010;
12'b10011111001010: data = 6'b111111;
12'b10011111001011: data = 6'b111111;
12'b10011111001100: data = 6'b111111;
12'b10011111001101: data = 6'b111111;
12'b10011111001110: data = 6'b111111;
12'b10011111001111: data = 6'b111111;
12'b10011111010000: data = 6'b111111;
12'b10011111010001: data = 6'b111111;
12'b10011111010010: data = 6'b111111;
12'b10011111010011: data = 6'b111111;
12'b10011111010100: data = 6'b111111;
12'b10011111010101: data = 6'b111111;
12'b10011111010110: data = 6'b111111;
12'b10011111010111: data = 6'b111111;
12'b10011111011000: data = 6'b111111;
12'b10011111011001: data = 6'b111111;
12'b10011111011010: data = 6'b111111;
12'b10011111011011: data = 6'b111111;
12'b10011111011100: data = 6'b111111;
12'b10011111011101: data = 6'b111111;
12'b10011111011110: data = 6'b111111;
12'b10011111011111: data = 6'b111111;
12'b10011111100000: data = 6'b111111;
12'b10011111100001: data = 6'b101010;
12'b10011111100010: data = 6'b010101;
12'b10011111100011: data = 6'b101001;
12'b10011111100100: data = 6'b101010;
12'b10011111100101: data = 6'b101010;
12'b10011111100110: data = 6'b101010;
12'b10011111100111: data = 6'b101010;
12'b10011111101000: data = 6'b101010;
12'b10011111101001: data = 6'b111111;
12'b10011111101010: data = 6'b111111;
12'b10011111101011: data = 6'b111111;
12'b10011111101100: data = 6'b111111;
12'b10011111101101: data = 6'b111111;
12'b10011111101110: data = 6'b111111;
12'b10011111101111: data = 6'b111111;
12'b10011111110000: data = 6'b111111;
12'b10011111110001: data = 6'b111111;
12'b10011111110010: data = 6'b111111;
12'b10011111110011: data = 6'b111111;
12'b10011111110100: data = 6'b111111;
12'b10011111110101: data = 6'b111111;
12'b10011111110110: data = 6'b111111;
12'b10011111110111: data = 6'b111111;
12'b10011111111000: data = 6'b111111;
12'b10011111111001: data = 6'b111111;
12'b10011111111010: data = 6'b111111;
12'b10011111111011: data = 6'b111111;
12'b10011111111100: data = 6'b111111;
12'b10011111111101: data = 6'b111111;
12'b10011111111110: data = 6'b111111;
12'b10011111111111: data = 6'b111111;
12'b100111110000000: data = 6'b111111;
12'b100111110000001: data = 6'b111111;
12'b100111110000010: data = 6'b111111;
12'b100111110000011: data = 6'b111111;
12'b100111110000100: data = 6'b101010;
12'b100111110000101: data = 6'b101010;
12'b100111110000110: data = 6'b101010;
12'b100111110000111: data = 6'b101010;
12'b100111110001000: data = 6'b101010;
12'b100111110001001: data = 6'b010101;
12'b100111110001010: data = 6'b010101;
12'b100111110001011: data = 6'b010101;
12'b100111110001100: data = 6'b000000;
12'b100111110001101: data = 6'b000000;
12'b100111110001110: data = 6'b101010;
12'b100111110001111: data = 6'b101010;
12'b100111110010000: data = 6'b101010;
12'b100111110010001: data = 6'b101010;
12'b100111110010010: data = 6'b010101;
12'b100111110010011: data = 6'b010101;
12'b100111110010100: data = 6'b010101;
12'b100111110010101: data = 6'b010101;
12'b100111110010110: data = 6'b010101;
12'b100111110010111: data = 6'b010101;
12'b100111110011000: data = 6'b010101;
12'b100111110011001: data = 6'b010101;
12'b100111110011010: data = 6'b010101;
12'b100111110011011: data = 6'b010101;
12'b100111110011100: data = 6'b010101;
12'b100111110011101: data = 6'b010101;
12'b100111110011110: data = 6'b010101;
12'b100111110011111: data = 6'b010101;
12'b100111110100000: data = 6'b010101;
12'b100111110100001: data = 6'b010101;
12'b100111110100010: data = 6'b010101;
12'b100111110100011: data = 6'b010101;
12'b100111110100100: data = 6'b010101;
12'b100111110100101: data = 6'b010101;
12'b100111110100110: data = 6'b010101;
12'b100111110100111: data = 6'b010101;
12'b100111110101000: data = 6'b010101;
12'b100111110101001: data = 6'b010101;
12'b100111110101010: data = 6'b010101;
12'b1010000000000: data = 6'b010101;
12'b1010000000001: data = 6'b010101;
12'b1010000000010: data = 6'b010101;
12'b1010000000011: data = 6'b010101;
12'b1010000000100: data = 6'b010101;
12'b1010000000101: data = 6'b010101;
12'b1010000000110: data = 6'b010101;
12'b1010000000111: data = 6'b010101;
12'b1010000001000: data = 6'b010101;
12'b1010000001001: data = 6'b010101;
12'b1010000001010: data = 6'b010101;
12'b1010000001011: data = 6'b010101;
12'b1010000001100: data = 6'b010101;
12'b1010000001101: data = 6'b010101;
12'b1010000001110: data = 6'b010101;
12'b1010000001111: data = 6'b010101;
12'b1010000010000: data = 6'b010101;
12'b1010000010001: data = 6'b010101;
12'b1010000010010: data = 6'b010101;
12'b1010000010011: data = 6'b010101;
12'b1010000010100: data = 6'b010101;
12'b1010000010101: data = 6'b010101;
12'b1010000010110: data = 6'b010101;
12'b1010000010111: data = 6'b010101;
12'b1010000011000: data = 6'b010101;
12'b1010000011001: data = 6'b101010;
12'b1010000011010: data = 6'b101010;
12'b1010000011011: data = 6'b101010;
12'b1010000011100: data = 6'b010101;
12'b1010000011101: data = 6'b000000;
12'b1010000011110: data = 6'b000000;
12'b1010000011111: data = 6'b010101;
12'b1010000100000: data = 6'b010101;
12'b1010000100001: data = 6'b010101;
12'b1010000100010: data = 6'b101010;
12'b1010000100011: data = 6'b101010;
12'b1010000100100: data = 6'b101010;
12'b1010000100101: data = 6'b101010;
12'b1010000100110: data = 6'b101010;
12'b1010000100111: data = 6'b101010;
12'b1010000101000: data = 6'b111111;
12'b1010000101001: data = 6'b111111;
12'b1010000101010: data = 6'b101010;
12'b1010000101011: data = 6'b101010;
12'b1010000101100: data = 6'b101010;
12'b1010000101101: data = 6'b101010;
12'b1010000101110: data = 6'b101010;
12'b1010000101111: data = 6'b101010;
12'b1010000110000: data = 6'b101010;
12'b1010000110001: data = 6'b101010;
12'b1010000110010: data = 6'b101010;
12'b1010000110011: data = 6'b101010;
12'b1010000110100: data = 6'b101010;
12'b1010000110101: data = 6'b101010;
12'b1010000110110: data = 6'b101010;
12'b1010000110111: data = 6'b101010;
12'b1010000111000: data = 6'b101010;
12'b1010000111001: data = 6'b101010;
12'b1010000111010: data = 6'b101010;
12'b1010000111011: data = 6'b101010;
12'b1010000111100: data = 6'b101010;
12'b1010000111101: data = 6'b101010;
12'b1010000111110: data = 6'b101010;
12'b1010000111111: data = 6'b111111;
12'b10100001000000: data = 6'b111111;
12'b10100001000001: data = 6'b101010;
12'b10100001000010: data = 6'b101010;
12'b10100001000011: data = 6'b101010;
12'b10100001000100: data = 6'b101010;
12'b10100001000101: data = 6'b101010;
12'b10100001000110: data = 6'b101010;
12'b10100001000111: data = 6'b101010;
12'b10100001001000: data = 6'b010101;
12'b10100001001001: data = 6'b101010;
12'b10100001001010: data = 6'b101010;
12'b10100001001011: data = 6'b101010;
12'b10100001001100: data = 6'b101010;
12'b10100001001101: data = 6'b101010;
12'b10100001001110: data = 6'b101010;
12'b10100001001111: data = 6'b101010;
12'b10100001010000: data = 6'b101010;
12'b10100001010001: data = 6'b101010;
12'b10100001010010: data = 6'b101010;
12'b10100001010011: data = 6'b101010;
12'b10100001010100: data = 6'b101010;
12'b10100001010101: data = 6'b101010;
12'b10100001010110: data = 6'b101010;
12'b10100001010111: data = 6'b101010;
12'b10100001011000: data = 6'b101010;
12'b10100001011001: data = 6'b101010;
12'b10100001011010: data = 6'b101010;
12'b10100001011011: data = 6'b101010;
12'b10100001011100: data = 6'b101010;
12'b10100001011101: data = 6'b101010;
12'b10100001011110: data = 6'b101010;
12'b10100001011111: data = 6'b101010;
12'b10100001100000: data = 6'b101010;
12'b10100001100001: data = 6'b101010;
12'b10100001100010: data = 6'b010101;
12'b10100001100011: data = 6'b101001;
12'b10100001100100: data = 6'b101010;
12'b10100001100101: data = 6'b101010;
12'b10100001100110: data = 6'b101010;
12'b10100001100111: data = 6'b101010;
12'b10100001101000: data = 6'b101010;
12'b10100001101001: data = 6'b101010;
12'b10100001101010: data = 6'b111111;
12'b10100001101011: data = 6'b101010;
12'b10100001101100: data = 6'b101010;
12'b10100001101101: data = 6'b101010;
12'b10100001101110: data = 6'b101010;
12'b10100001101111: data = 6'b101010;
12'b10100001110000: data = 6'b101010;
12'b10100001110001: data = 6'b101010;
12'b10100001110010: data = 6'b111111;
12'b10100001110011: data = 6'b101010;
12'b10100001110100: data = 6'b101010;
12'b10100001110101: data = 6'b101010;
12'b10100001110110: data = 6'b101010;
12'b10100001110111: data = 6'b101010;
12'b10100001111000: data = 6'b101010;
12'b10100001111001: data = 6'b101010;
12'b10100001111010: data = 6'b101010;
12'b10100001111011: data = 6'b101010;
12'b10100001111100: data = 6'b101010;
12'b10100001111101: data = 6'b101010;
12'b10100001111110: data = 6'b101010;
12'b10100001111111: data = 6'b101010;
12'b101000010000000: data = 6'b101010;
12'b101000010000001: data = 6'b101010;
12'b101000010000010: data = 6'b101010;
12'b101000010000011: data = 6'b101010;
12'b101000010000100: data = 6'b101010;
12'b101000010000101: data = 6'b101010;
12'b101000010000110: data = 6'b101010;
12'b101000010000111: data = 6'b101010;
12'b101000010001000: data = 6'b101010;
12'b101000010001001: data = 6'b010101;
12'b101000010001010: data = 6'b010101;
12'b101000010001011: data = 6'b010101;
12'b101000010001100: data = 6'b000000;
12'b101000010001101: data = 6'b000000;
12'b101000010001110: data = 6'b101010;
12'b101000010001111: data = 6'b101010;
12'b101000010010000: data = 6'b101010;
12'b101000010010001: data = 6'b101010;
12'b101000010010010: data = 6'b010101;
12'b101000010010011: data = 6'b010101;
12'b101000010010100: data = 6'b010101;
12'b101000010010101: data = 6'b010101;
12'b101000010010110: data = 6'b010101;
12'b101000010010111: data = 6'b010101;
12'b101000010011000: data = 6'b010101;
12'b101000010011001: data = 6'b010101;
12'b101000010011010: data = 6'b010101;
12'b101000010011011: data = 6'b010101;
12'b101000010011100: data = 6'b010101;
12'b101000010011101: data = 6'b010101;
12'b101000010011110: data = 6'b010101;
12'b101000010011111: data = 6'b010101;
12'b101000010100000: data = 6'b010101;
12'b101000010100001: data = 6'b010101;
12'b101000010100010: data = 6'b010101;
12'b101000010100011: data = 6'b010101;
12'b101000010100100: data = 6'b010101;
12'b101000010100101: data = 6'b010101;
12'b101000010100110: data = 6'b010101;
12'b101000010100111: data = 6'b010101;
12'b101000010101000: data = 6'b010101;
12'b101000010101001: data = 6'b010101;
12'b101000010101010: data = 6'b010101;
12'b1010001000000: data = 6'b010101;
12'b1010001000001: data = 6'b010101;
12'b1010001000010: data = 6'b010101;
12'b1010001000011: data = 6'b010101;
12'b1010001000100: data = 6'b010101;
12'b1010001000101: data = 6'b010101;
12'b1010001000110: data = 6'b010101;
12'b1010001000111: data = 6'b010101;
12'b1010001001000: data = 6'b010101;
12'b1010001001001: data = 6'b010101;
12'b1010001001010: data = 6'b010101;
12'b1010001001011: data = 6'b010101;
12'b1010001001100: data = 6'b010101;
12'b1010001001101: data = 6'b010101;
12'b1010001001110: data = 6'b010101;
12'b1010001001111: data = 6'b010101;
12'b1010001010000: data = 6'b010101;
12'b1010001010001: data = 6'b010101;
12'b1010001010010: data = 6'b010101;
12'b1010001010011: data = 6'b010101;
12'b1010001010100: data = 6'b010101;
12'b1010001010101: data = 6'b010101;
12'b1010001010110: data = 6'b010101;
12'b1010001010111: data = 6'b010101;
12'b1010001011000: data = 6'b010101;
12'b1010001011001: data = 6'b101010;
12'b1010001011010: data = 6'b101010;
12'b1010001011011: data = 6'b101010;
12'b1010001011100: data = 6'b010101;
12'b1010001011101: data = 6'b000000;
12'b1010001011110: data = 6'b000000;
12'b1010001011111: data = 6'b010101;
12'b1010001100000: data = 6'b010101;
12'b1010001100001: data = 6'b010101;
12'b1010001100010: data = 6'b101010;
12'b1010001100011: data = 6'b101010;
12'b1010001100100: data = 6'b101010;
12'b1010001100101: data = 6'b101010;
12'b1010001100110: data = 6'b101010;
12'b1010001100111: data = 6'b101010;
12'b1010001101000: data = 6'b101010;
12'b1010001101001: data = 6'b101010;
12'b1010001101010: data = 6'b101010;
12'b1010001101011: data = 6'b101010;
12'b1010001101100: data = 6'b101010;
12'b1010001101101: data = 6'b101010;
12'b1010001101110: data = 6'b101010;
12'b1010001101111: data = 6'b101010;
12'b1010001110000: data = 6'b101010;
12'b1010001110001: data = 6'b101010;
12'b1010001110010: data = 6'b101010;
12'b1010001110011: data = 6'b101010;
12'b1010001110100: data = 6'b101010;
12'b1010001110101: data = 6'b101010;
12'b1010001110110: data = 6'b101010;
12'b1010001110111: data = 6'b101010;
12'b1010001111000: data = 6'b101010;
12'b1010001111001: data = 6'b101010;
12'b1010001111010: data = 6'b101010;
12'b1010001111011: data = 6'b101010;
12'b1010001111100: data = 6'b101010;
12'b1010001111101: data = 6'b101010;
12'b1010001111110: data = 6'b101010;
12'b1010001111111: data = 6'b101010;
12'b10100011000000: data = 6'b101010;
12'b10100011000001: data = 6'b101010;
12'b10100011000010: data = 6'b101010;
12'b10100011000011: data = 6'b101010;
12'b10100011000100: data = 6'b101010;
12'b10100011000101: data = 6'b101010;
12'b10100011000110: data = 6'b101010;
12'b10100011000111: data = 6'b101010;
12'b10100011001000: data = 6'b101001;
12'b10100011001001: data = 6'b101010;
12'b10100011001010: data = 6'b101010;
12'b10100011001011: data = 6'b101010;
12'b10100011001100: data = 6'b101010;
12'b10100011001101: data = 6'b101010;
12'b10100011001110: data = 6'b101010;
12'b10100011001111: data = 6'b101010;
12'b10100011010000: data = 6'b101010;
12'b10100011010001: data = 6'b101010;
12'b10100011010010: data = 6'b101010;
12'b10100011010011: data = 6'b101010;
12'b10100011010100: data = 6'b101010;
12'b10100011010101: data = 6'b101010;
12'b10100011010110: data = 6'b101010;
12'b10100011010111: data = 6'b101010;
12'b10100011011000: data = 6'b101010;
12'b10100011011001: data = 6'b101010;
12'b10100011011010: data = 6'b101010;
12'b10100011011011: data = 6'b101010;
12'b10100011011100: data = 6'b101010;
12'b10100011011101: data = 6'b101010;
12'b10100011011110: data = 6'b101010;
12'b10100011011111: data = 6'b101010;
12'b10100011100000: data = 6'b101010;
12'b10100011100001: data = 6'b101010;
12'b10100011100010: data = 6'b010101;
12'b10100011100011: data = 6'b101001;
12'b10100011100100: data = 6'b101010;
12'b10100011100101: data = 6'b101010;
12'b10100011100110: data = 6'b101010;
12'b10100011100111: data = 6'b101010;
12'b10100011101000: data = 6'b101010;
12'b10100011101001: data = 6'b101010;
12'b10100011101010: data = 6'b101010;
12'b10100011101011: data = 6'b101010;
12'b10100011101100: data = 6'b101010;
12'b10100011101101: data = 6'b101010;
12'b10100011101110: data = 6'b101010;
12'b10100011101111: data = 6'b101010;
12'b10100011110000: data = 6'b101010;
12'b10100011110001: data = 6'b101010;
12'b10100011110010: data = 6'b101010;
12'b10100011110011: data = 6'b101010;
12'b10100011110100: data = 6'b101010;
12'b10100011110101: data = 6'b101010;
12'b10100011110110: data = 6'b101010;
12'b10100011110111: data = 6'b101010;
12'b10100011111000: data = 6'b101010;
12'b10100011111001: data = 6'b101010;
12'b10100011111010: data = 6'b101010;
12'b10100011111011: data = 6'b101010;
12'b10100011111100: data = 6'b101010;
12'b10100011111101: data = 6'b101010;
12'b10100011111110: data = 6'b101010;
12'b10100011111111: data = 6'b101010;
12'b101000110000000: data = 6'b101010;
12'b101000110000001: data = 6'b101010;
12'b101000110000010: data = 6'b101010;
12'b101000110000011: data = 6'b101010;
12'b101000110000100: data = 6'b101010;
12'b101000110000101: data = 6'b101010;
12'b101000110000110: data = 6'b101010;
12'b101000110000111: data = 6'b101010;
12'b101000110001000: data = 6'b101010;
12'b101000110001001: data = 6'b010101;
12'b101000110001010: data = 6'b010101;
12'b101000110001011: data = 6'b010101;
12'b101000110001100: data = 6'b000000;
12'b101000110001101: data = 6'b000000;
12'b101000110001110: data = 6'b101010;
12'b101000110001111: data = 6'b101010;
12'b101000110010000: data = 6'b101010;
12'b101000110010001: data = 6'b101010;
12'b101000110010010: data = 6'b010101;
12'b101000110010011: data = 6'b010101;
12'b101000110010100: data = 6'b010101;
12'b101000110010101: data = 6'b010101;
12'b101000110010110: data = 6'b010101;
12'b101000110010111: data = 6'b010101;
12'b101000110011000: data = 6'b010101;
12'b101000110011001: data = 6'b010101;
12'b101000110011010: data = 6'b010101;
12'b101000110011011: data = 6'b010101;
12'b101000110011100: data = 6'b010101;
12'b101000110011101: data = 6'b010101;
12'b101000110011110: data = 6'b010101;
12'b101000110011111: data = 6'b010101;
12'b101000110100000: data = 6'b010101;
12'b101000110100001: data = 6'b010101;
12'b101000110100010: data = 6'b010101;
12'b101000110100011: data = 6'b010101;
12'b101000110100100: data = 6'b010101;
12'b101000110100101: data = 6'b010101;
12'b101000110100110: data = 6'b010101;
12'b101000110100111: data = 6'b010101;
12'b101000110101000: data = 6'b010101;
12'b101000110101001: data = 6'b010101;
12'b101000110101010: data = 6'b010101;
12'b1010010000000: data = 6'b010101;
12'b1010010000001: data = 6'b010101;
12'b1010010000010: data = 6'b010101;
12'b1010010000011: data = 6'b010101;
12'b1010010000100: data = 6'b010101;
12'b1010010000101: data = 6'b010101;
12'b1010010000110: data = 6'b010101;
12'b1010010000111: data = 6'b010101;
12'b1010010001000: data = 6'b010101;
12'b1010010001001: data = 6'b010101;
12'b1010010001010: data = 6'b010101;
12'b1010010001011: data = 6'b010101;
12'b1010010001100: data = 6'b010101;
12'b1010010001101: data = 6'b010101;
12'b1010010001110: data = 6'b010101;
12'b1010010001111: data = 6'b010101;
12'b1010010010000: data = 6'b010101;
12'b1010010010001: data = 6'b010101;
12'b1010010010010: data = 6'b010101;
12'b1010010010011: data = 6'b010101;
12'b1010010010100: data = 6'b010101;
12'b1010010010101: data = 6'b010101;
12'b1010010010110: data = 6'b010101;
12'b1010010010111: data = 6'b010101;
12'b1010010011000: data = 6'b010101;
12'b1010010011001: data = 6'b101010;
12'b1010010011010: data = 6'b101010;
12'b1010010011011: data = 6'b101010;
12'b1010010011100: data = 6'b010101;
12'b1010010011101: data = 6'b000000;
12'b1010010011110: data = 6'b000000;
12'b1010010011111: data = 6'b010101;
12'b1010010100000: data = 6'b010101;
12'b1010010100001: data = 6'b010101;
12'b1010010100010: data = 6'b101010;
12'b1010010100011: data = 6'b101010;
12'b1010010100100: data = 6'b101010;
12'b1010010100101: data = 6'b101010;
12'b1010010100110: data = 6'b101010;
12'b1010010100111: data = 6'b101010;
12'b1010010101000: data = 6'b101010;
12'b1010010101001: data = 6'b101010;
12'b1010010101010: data = 6'b101010;
12'b1010010101011: data = 6'b101010;
12'b1010010101100: data = 6'b101010;
12'b1010010101101: data = 6'b101010;
12'b1010010101110: data = 6'b101010;
12'b1010010101111: data = 6'b101010;
12'b1010010110000: data = 6'b101010;
12'b1010010110001: data = 6'b101010;
12'b1010010110010: data = 6'b101010;
12'b1010010110011: data = 6'b101010;
12'b1010010110100: data = 6'b101010;
12'b1010010110101: data = 6'b101010;
12'b1010010110110: data = 6'b101010;
12'b1010010110111: data = 6'b101010;
12'b1010010111000: data = 6'b101010;
12'b1010010111001: data = 6'b101010;
12'b1010010111010: data = 6'b101010;
12'b1010010111011: data = 6'b101010;
12'b1010010111100: data = 6'b101010;
12'b1010010111101: data = 6'b101010;
12'b1010010111110: data = 6'b101010;
12'b1010010111111: data = 6'b101010;
12'b10100101000000: data = 6'b101010;
12'b10100101000001: data = 6'b101010;
12'b10100101000010: data = 6'b101010;
12'b10100101000011: data = 6'b101010;
12'b10100101000100: data = 6'b101010;
12'b10100101000101: data = 6'b101010;
12'b10100101000110: data = 6'b101010;
12'b10100101000111: data = 6'b101010;
12'b10100101001000: data = 6'b101001;
12'b10100101001001: data = 6'b101010;
12'b10100101001010: data = 6'b101010;
12'b10100101001011: data = 6'b101010;
12'b10100101001100: data = 6'b101010;
12'b10100101001101: data = 6'b101010;
12'b10100101001110: data = 6'b101010;
12'b10100101001111: data = 6'b101010;
12'b10100101010000: data = 6'b101010;
12'b10100101010001: data = 6'b101010;
12'b10100101010010: data = 6'b101010;
12'b10100101010011: data = 6'b101010;
12'b10100101010100: data = 6'b101010;
12'b10100101010101: data = 6'b101010;
12'b10100101010110: data = 6'b101010;
12'b10100101010111: data = 6'b101010;
12'b10100101011000: data = 6'b101010;
12'b10100101011001: data = 6'b101010;
12'b10100101011010: data = 6'b101010;
12'b10100101011011: data = 6'b101010;
12'b10100101011100: data = 6'b101010;
12'b10100101011101: data = 6'b101010;
12'b10100101011110: data = 6'b101010;
12'b10100101011111: data = 6'b101010;
12'b10100101100000: data = 6'b101010;
12'b10100101100001: data = 6'b101010;
12'b10100101100010: data = 6'b010101;
12'b10100101100011: data = 6'b101001;
12'b10100101100100: data = 6'b101010;
12'b10100101100101: data = 6'b101010;
12'b10100101100110: data = 6'b101010;
12'b10100101100111: data = 6'b101010;
12'b10100101101000: data = 6'b101010;
12'b10100101101001: data = 6'b101010;
12'b10100101101010: data = 6'b101010;
12'b10100101101011: data = 6'b101010;
12'b10100101101100: data = 6'b101010;
12'b10100101101101: data = 6'b101010;
12'b10100101101110: data = 6'b101010;
12'b10100101101111: data = 6'b101010;
12'b10100101110000: data = 6'b101010;
12'b10100101110001: data = 6'b101010;
12'b10100101110010: data = 6'b101010;
12'b10100101110011: data = 6'b101010;
12'b10100101110100: data = 6'b101010;
12'b10100101110101: data = 6'b101010;
12'b10100101110110: data = 6'b101010;
12'b10100101110111: data = 6'b101010;
12'b10100101111000: data = 6'b101010;
12'b10100101111001: data = 6'b101010;
12'b10100101111010: data = 6'b101010;
12'b10100101111011: data = 6'b101010;
12'b10100101111100: data = 6'b101010;
12'b10100101111101: data = 6'b101010;
12'b10100101111110: data = 6'b101010;
12'b10100101111111: data = 6'b101010;
12'b101001010000000: data = 6'b101010;
12'b101001010000001: data = 6'b101010;
12'b101001010000010: data = 6'b101010;
12'b101001010000011: data = 6'b101010;
12'b101001010000100: data = 6'b101010;
12'b101001010000101: data = 6'b101010;
12'b101001010000110: data = 6'b101010;
12'b101001010000111: data = 6'b101010;
12'b101001010001000: data = 6'b101010;
12'b101001010001001: data = 6'b010101;
12'b101001010001010: data = 6'b010101;
12'b101001010001011: data = 6'b010101;
12'b101001010001100: data = 6'b000000;
12'b101001010001101: data = 6'b000000;
12'b101001010001110: data = 6'b101010;
12'b101001010001111: data = 6'b101010;
12'b101001010010000: data = 6'b101010;
12'b101001010010001: data = 6'b101010;
12'b101001010010010: data = 6'b010101;
12'b101001010010011: data = 6'b010101;
12'b101001010010100: data = 6'b010101;
12'b101001010010101: data = 6'b010101;
12'b101001010010110: data = 6'b010101;
12'b101001010010111: data = 6'b010101;
12'b101001010011000: data = 6'b010101;
12'b101001010011001: data = 6'b010101;
12'b101001010011010: data = 6'b010101;
12'b101001010011011: data = 6'b010101;
12'b101001010011100: data = 6'b010101;
12'b101001010011101: data = 6'b010101;
12'b101001010011110: data = 6'b010101;
12'b101001010011111: data = 6'b010101;
12'b101001010100000: data = 6'b010101;
12'b101001010100001: data = 6'b010101;
12'b101001010100010: data = 6'b010101;
12'b101001010100011: data = 6'b010101;
12'b101001010100100: data = 6'b010101;
12'b101001010100101: data = 6'b010101;
12'b101001010100110: data = 6'b010101;
12'b101001010100111: data = 6'b010101;
12'b101001010101000: data = 6'b010101;
12'b101001010101001: data = 6'b010101;
12'b101001010101010: data = 6'b010101;
12'b1010011000000: data = 6'b010101;
12'b1010011000001: data = 6'b010101;
12'b1010011000010: data = 6'b010101;
12'b1010011000011: data = 6'b010101;
12'b1010011000100: data = 6'b010101;
12'b1010011000101: data = 6'b010101;
12'b1010011000110: data = 6'b010101;
12'b1010011000111: data = 6'b010101;
12'b1010011001000: data = 6'b010101;
12'b1010011001001: data = 6'b010101;
12'b1010011001010: data = 6'b010101;
12'b1010011001011: data = 6'b010101;
12'b1010011001100: data = 6'b010101;
12'b1010011001101: data = 6'b010101;
12'b1010011001110: data = 6'b010101;
12'b1010011001111: data = 6'b010101;
12'b1010011010000: data = 6'b010101;
12'b1010011010001: data = 6'b010101;
12'b1010011010010: data = 6'b010101;
12'b1010011010011: data = 6'b010101;
12'b1010011010100: data = 6'b010101;
12'b1010011010101: data = 6'b010101;
12'b1010011010110: data = 6'b010101;
12'b1010011010111: data = 6'b010101;
12'b1010011011000: data = 6'b010101;
12'b1010011011001: data = 6'b101010;
12'b1010011011010: data = 6'b101010;
12'b1010011011011: data = 6'b101010;
12'b1010011011100: data = 6'b010101;
12'b1010011011101: data = 6'b000000;
12'b1010011011110: data = 6'b000000;
12'b1010011011111: data = 6'b010101;
12'b1010011100000: data = 6'b010101;
12'b1010011100001: data = 6'b010101;
12'b1010011100010: data = 6'b101010;
12'b1010011100011: data = 6'b101010;
12'b1010011100100: data = 6'b101010;
12'b1010011100101: data = 6'b101010;
12'b1010011100110: data = 6'b101010;
12'b1010011100111: data = 6'b101010;
12'b1010011101000: data = 6'b101001;
12'b1010011101001: data = 6'b101001;
12'b1010011101010: data = 6'b101010;
12'b1010011101011: data = 6'b101010;
12'b1010011101100: data = 6'b101010;
12'b1010011101101: data = 6'b101010;
12'b1010011101110: data = 6'b101010;
12'b1010011101111: data = 6'b101010;
12'b1010011110000: data = 6'b101010;
12'b1010011110001: data = 6'b101010;
12'b1010011110010: data = 6'b101010;
12'b1010011110011: data = 6'b101010;
12'b1010011110100: data = 6'b101010;
12'b1010011110101: data = 6'b101010;
12'b1010011110110: data = 6'b101010;
12'b1010011110111: data = 6'b101010;
12'b1010011111000: data = 6'b101010;
12'b1010011111001: data = 6'b101010;
12'b1010011111010: data = 6'b101010;
12'b1010011111011: data = 6'b101010;
12'b1010011111100: data = 6'b101010;
12'b1010011111101: data = 6'b101010;
12'b1010011111110: data = 6'b101010;
12'b1010011111111: data = 6'b101010;
12'b10100111000000: data = 6'b101010;
12'b10100111000001: data = 6'b101010;
12'b10100111000010: data = 6'b101010;
12'b10100111000011: data = 6'b101010;
12'b10100111000100: data = 6'b101010;
12'b10100111000101: data = 6'b101010;
12'b10100111000110: data = 6'b101010;
12'b10100111000111: data = 6'b101010;
12'b10100111001000: data = 6'b101010;
12'b10100111001001: data = 6'b101010;
12'b10100111001010: data = 6'b101010;
12'b10100111001011: data = 6'b101010;
12'b10100111001100: data = 6'b101010;
12'b10100111001101: data = 6'b101010;
12'b10100111001110: data = 6'b101010;
12'b10100111001111: data = 6'b101010;
12'b10100111010000: data = 6'b101010;
12'b10100111010001: data = 6'b101010;
12'b10100111010010: data = 6'b101010;
12'b10100111010011: data = 6'b101010;
12'b10100111010100: data = 6'b101010;
12'b10100111010101: data = 6'b101010;
12'b10100111010110: data = 6'b101010;
12'b10100111010111: data = 6'b101010;
12'b10100111011000: data = 6'b101010;
12'b10100111011001: data = 6'b101010;
12'b10100111011010: data = 6'b101010;
12'b10100111011011: data = 6'b101010;
12'b10100111011100: data = 6'b101010;
12'b10100111011101: data = 6'b101010;
12'b10100111011110: data = 6'b101010;
12'b10100111011111: data = 6'b101010;
12'b10100111100000: data = 6'b101010;
12'b10100111100001: data = 6'b101001;
12'b10100111100010: data = 6'b010101;
12'b10100111100011: data = 6'b101001;
12'b10100111100100: data = 6'b101010;
12'b10100111100101: data = 6'b101010;
12'b10100111100110: data = 6'b101010;
12'b10100111100111: data = 6'b101010;
12'b10100111101000: data = 6'b101010;
12'b10100111101001: data = 6'b101010;
12'b10100111101010: data = 6'b101010;
12'b10100111101011: data = 6'b101010;
12'b10100111101100: data = 6'b101010;
12'b10100111101101: data = 6'b101010;
12'b10100111101110: data = 6'b101010;
12'b10100111101111: data = 6'b101010;
12'b10100111110000: data = 6'b101010;
12'b10100111110001: data = 6'b101010;
12'b10100111110010: data = 6'b101010;
12'b10100111110011: data = 6'b101010;
12'b10100111110100: data = 6'b101010;
12'b10100111110101: data = 6'b101010;
12'b10100111110110: data = 6'b101010;
12'b10100111110111: data = 6'b101010;
12'b10100111111000: data = 6'b101010;
12'b10100111111001: data = 6'b101010;
12'b10100111111010: data = 6'b101010;
12'b10100111111011: data = 6'b101010;
12'b10100111111100: data = 6'b101010;
12'b10100111111101: data = 6'b101010;
12'b10100111111110: data = 6'b101010;
12'b10100111111111: data = 6'b101010;
12'b101001110000000: data = 6'b101010;
12'b101001110000001: data = 6'b101010;
12'b101001110000010: data = 6'b101010;
12'b101001110000011: data = 6'b101010;
12'b101001110000100: data = 6'b101010;
12'b101001110000101: data = 6'b101010;
12'b101001110000110: data = 6'b101010;
12'b101001110000111: data = 6'b101010;
12'b101001110001000: data = 6'b101010;
12'b101001110001001: data = 6'b010101;
12'b101001110001010: data = 6'b010101;
12'b101001110001011: data = 6'b010101;
12'b101001110001100: data = 6'b000000;
12'b101001110001101: data = 6'b000000;
12'b101001110001110: data = 6'b101010;
12'b101001110001111: data = 6'b101010;
12'b101001110010000: data = 6'b101010;
12'b101001110010001: data = 6'b101010;
12'b101001110010010: data = 6'b010101;
12'b101001110010011: data = 6'b010101;
12'b101001110010100: data = 6'b010101;
12'b101001110010101: data = 6'b010101;
12'b101001110010110: data = 6'b010101;
12'b101001110010111: data = 6'b010101;
12'b101001110011000: data = 6'b010101;
12'b101001110011001: data = 6'b010101;
12'b101001110011010: data = 6'b010101;
12'b101001110011011: data = 6'b010101;
12'b101001110011100: data = 6'b010101;
12'b101001110011101: data = 6'b010101;
12'b101001110011110: data = 6'b010101;
12'b101001110011111: data = 6'b010101;
12'b101001110100000: data = 6'b010101;
12'b101001110100001: data = 6'b010101;
12'b101001110100010: data = 6'b010101;
12'b101001110100011: data = 6'b010101;
12'b101001110100100: data = 6'b010101;
12'b101001110100101: data = 6'b010101;
12'b101001110100110: data = 6'b010101;
12'b101001110100111: data = 6'b010101;
12'b101001110101000: data = 6'b010101;
12'b101001110101001: data = 6'b010101;
12'b101001110101010: data = 6'b010101;
12'b1010100000000: data = 6'b010101;
12'b1010100000001: data = 6'b010101;
12'b1010100000010: data = 6'b010101;
12'b1010100000011: data = 6'b010101;
12'b1010100000100: data = 6'b010101;
12'b1010100000101: data = 6'b010101;
12'b1010100000110: data = 6'b010101;
12'b1010100000111: data = 6'b010101;
12'b1010100001000: data = 6'b010101;
12'b1010100001001: data = 6'b010101;
12'b1010100001010: data = 6'b010101;
12'b1010100001011: data = 6'b010101;
12'b1010100001100: data = 6'b010101;
12'b1010100001101: data = 6'b010101;
12'b1010100001110: data = 6'b010101;
12'b1010100001111: data = 6'b010101;
12'b1010100010000: data = 6'b010101;
12'b1010100010001: data = 6'b010101;
12'b1010100010010: data = 6'b010101;
12'b1010100010011: data = 6'b010101;
12'b1010100010100: data = 6'b010101;
12'b1010100010101: data = 6'b010101;
12'b1010100010110: data = 6'b010101;
12'b1010100010111: data = 6'b010101;
12'b1010100011000: data = 6'b010101;
12'b1010100011001: data = 6'b101010;
12'b1010100011010: data = 6'b101010;
12'b1010100011011: data = 6'b101010;
12'b1010100011100: data = 6'b010101;
12'b1010100011101: data = 6'b000000;
12'b1010100011110: data = 6'b000000;
12'b1010100011111: data = 6'b010101;
12'b1010100100000: data = 6'b010101;
12'b1010100100001: data = 6'b010101;
12'b1010100100010: data = 6'b101010;
12'b1010100100011: data = 6'b101010;
12'b1010100100100: data = 6'b101010;
12'b1010100100101: data = 6'b101010;
12'b1010100100110: data = 6'b101010;
12'b1010100100111: data = 6'b101010;
12'b1010100101000: data = 6'b101001;
12'b1010100101001: data = 6'b101001;
12'b1010100101010: data = 6'b101010;
12'b1010100101011: data = 6'b101010;
12'b1010100101100: data = 6'b101010;
12'b1010100101101: data = 6'b101010;
12'b1010100101110: data = 6'b101010;
12'b1010100101111: data = 6'b101010;
12'b1010100110000: data = 6'b101010;
12'b1010100110001: data = 6'b101010;
12'b1010100110010: data = 6'b101010;
12'b1010100110011: data = 6'b101010;
12'b1010100110100: data = 6'b101010;
12'b1010100110101: data = 6'b101010;
12'b1010100110110: data = 6'b101010;
12'b1010100110111: data = 6'b101010;
12'b1010100111000: data = 6'b101010;
12'b1010100111001: data = 6'b101010;
12'b1010100111010: data = 6'b101010;
12'b1010100111011: data = 6'b101010;
12'b1010100111100: data = 6'b101010;
12'b1010100111101: data = 6'b101010;
12'b1010100111110: data = 6'b101010;
12'b1010100111111: data = 6'b101010;
12'b10101001000000: data = 6'b101010;
12'b10101001000001: data = 6'b101010;
12'b10101001000010: data = 6'b101010;
12'b10101001000011: data = 6'b101010;
12'b10101001000100: data = 6'b101010;
12'b10101001000101: data = 6'b101010;
12'b10101001000110: data = 6'b101010;
12'b10101001000111: data = 6'b101010;
12'b10101001001000: data = 6'b101010;
12'b10101001001001: data = 6'b101010;
12'b10101001001010: data = 6'b101010;
12'b10101001001011: data = 6'b101010;
12'b10101001001100: data = 6'b101010;
12'b10101001001101: data = 6'b101010;
12'b10101001001110: data = 6'b101010;
12'b10101001001111: data = 6'b101010;
12'b10101001010000: data = 6'b101010;
12'b10101001010001: data = 6'b101010;
12'b10101001010010: data = 6'b101010;
12'b10101001010011: data = 6'b101010;
12'b10101001010100: data = 6'b101010;
12'b10101001010101: data = 6'b101010;
12'b10101001010110: data = 6'b101010;
12'b10101001010111: data = 6'b101010;
12'b10101001011000: data = 6'b101010;
12'b10101001011001: data = 6'b101010;
12'b10101001011010: data = 6'b101010;
12'b10101001011011: data = 6'b101010;
12'b10101001011100: data = 6'b101010;
12'b10101001011101: data = 6'b101010;
12'b10101001011110: data = 6'b101010;
12'b10101001011111: data = 6'b101010;
12'b10101001100000: data = 6'b101010;
12'b10101001100001: data = 6'b101001;
12'b10101001100010: data = 6'b010101;
12'b10101001100011: data = 6'b101001;
12'b10101001100100: data = 6'b101010;
12'b10101001100101: data = 6'b101010;
12'b10101001100110: data = 6'b101010;
12'b10101001100111: data = 6'b101010;
12'b10101001101000: data = 6'b101010;
12'b10101001101001: data = 6'b101010;
12'b10101001101010: data = 6'b101010;
12'b10101001101011: data = 6'b101010;
12'b10101001101100: data = 6'b101010;
12'b10101001101101: data = 6'b101010;
12'b10101001101110: data = 6'b101010;
12'b10101001101111: data = 6'b101010;
12'b10101001110000: data = 6'b101010;
12'b10101001110001: data = 6'b101010;
12'b10101001110010: data = 6'b101010;
12'b10101001110011: data = 6'b101010;
12'b10101001110100: data = 6'b101010;
12'b10101001110101: data = 6'b101010;
12'b10101001110110: data = 6'b101010;
12'b10101001110111: data = 6'b101010;
12'b10101001111000: data = 6'b101010;
12'b10101001111001: data = 6'b101010;
12'b10101001111010: data = 6'b101010;
12'b10101001111011: data = 6'b101010;
12'b10101001111100: data = 6'b101010;
12'b10101001111101: data = 6'b101010;
12'b10101001111110: data = 6'b101010;
12'b10101001111111: data = 6'b101010;
12'b101010010000000: data = 6'b101010;
12'b101010010000001: data = 6'b101010;
12'b101010010000010: data = 6'b101010;
12'b101010010000011: data = 6'b101010;
12'b101010010000100: data = 6'b101010;
12'b101010010000101: data = 6'b101010;
12'b101010010000110: data = 6'b101010;
12'b101010010000111: data = 6'b101010;
12'b101010010001000: data = 6'b101010;
12'b101010010001001: data = 6'b010101;
12'b101010010001010: data = 6'b010101;
12'b101010010001011: data = 6'b010101;
12'b101010010001100: data = 6'b000000;
12'b101010010001101: data = 6'b000000;
12'b101010010001110: data = 6'b101010;
12'b101010010001111: data = 6'b101010;
12'b101010010010000: data = 6'b101010;
12'b101010010010001: data = 6'b101010;
12'b101010010010010: data = 6'b010101;
12'b101010010010011: data = 6'b010101;
12'b101010010010100: data = 6'b010101;
12'b101010010010101: data = 6'b010101;
12'b101010010010110: data = 6'b010101;
12'b101010010010111: data = 6'b010101;
12'b101010010011000: data = 6'b010101;
12'b101010010011001: data = 6'b010101;
12'b101010010011010: data = 6'b010101;
12'b101010010011011: data = 6'b010101;
12'b101010010011100: data = 6'b010101;
12'b101010010011101: data = 6'b010101;
12'b101010010011110: data = 6'b010101;
12'b101010010011111: data = 6'b010101;
12'b101010010100000: data = 6'b010101;
12'b101010010100001: data = 6'b010101;
12'b101010010100010: data = 6'b010101;
12'b101010010100011: data = 6'b010101;
12'b101010010100100: data = 6'b010101;
12'b101010010100101: data = 6'b010101;
12'b101010010100110: data = 6'b010101;
12'b101010010100111: data = 6'b010101;
12'b101010010101000: data = 6'b010101;
12'b101010010101001: data = 6'b010101;
12'b101010010101010: data = 6'b010101;
12'b1010101000000: data = 6'b010101;
12'b1010101000001: data = 6'b010101;
12'b1010101000010: data = 6'b010101;
12'b1010101000011: data = 6'b010101;
12'b1010101000100: data = 6'b010101;
12'b1010101000101: data = 6'b010101;
12'b1010101000110: data = 6'b010101;
12'b1010101000111: data = 6'b010101;
12'b1010101001000: data = 6'b010101;
12'b1010101001001: data = 6'b010101;
12'b1010101001010: data = 6'b010101;
12'b1010101001011: data = 6'b010101;
12'b1010101001100: data = 6'b010101;
12'b1010101001101: data = 6'b010101;
12'b1010101001110: data = 6'b010101;
12'b1010101001111: data = 6'b010101;
12'b1010101010000: data = 6'b010101;
12'b1010101010001: data = 6'b010101;
12'b1010101010010: data = 6'b010101;
12'b1010101010011: data = 6'b010101;
12'b1010101010100: data = 6'b010101;
12'b1010101010101: data = 6'b010101;
12'b1010101010110: data = 6'b010101;
12'b1010101010111: data = 6'b010101;
12'b1010101011000: data = 6'b010101;
12'b1010101011001: data = 6'b101010;
12'b1010101011010: data = 6'b101010;
12'b1010101011011: data = 6'b101010;
12'b1010101011100: data = 6'b010101;
12'b1010101011101: data = 6'b000000;
12'b1010101011110: data = 6'b000000;
12'b1010101011111: data = 6'b010101;
12'b1010101100000: data = 6'b010101;
12'b1010101100001: data = 6'b010101;
12'b1010101100010: data = 6'b101010;
12'b1010101100011: data = 6'b101010;
12'b1010101100100: data = 6'b101010;
12'b1010101100101: data = 6'b101010;
12'b1010101100110: data = 6'b101010;
12'b1010101100111: data = 6'b101010;
12'b1010101101000: data = 6'b101010;
12'b1010101101001: data = 6'b101010;
12'b1010101101010: data = 6'b101010;
12'b1010101101011: data = 6'b101010;
12'b1010101101100: data = 6'b101010;
12'b1010101101101: data = 6'b101010;
12'b1010101101110: data = 6'b101010;
12'b1010101101111: data = 6'b101010;
12'b1010101110000: data = 6'b101010;
12'b1010101110001: data = 6'b101010;
12'b1010101110010: data = 6'b101010;
12'b1010101110011: data = 6'b101010;
12'b1010101110100: data = 6'b101010;
12'b1010101110101: data = 6'b101010;
12'b1010101110110: data = 6'b101010;
12'b1010101110111: data = 6'b101010;
12'b1010101111000: data = 6'b101010;
12'b1010101111001: data = 6'b101010;
12'b1010101111010: data = 6'b101010;
12'b1010101111011: data = 6'b101010;
12'b1010101111100: data = 6'b101010;
12'b1010101111101: data = 6'b101010;
12'b1010101111110: data = 6'b101010;
12'b1010101111111: data = 6'b101010;
12'b10101011000000: data = 6'b101010;
12'b10101011000001: data = 6'b101010;
12'b10101011000010: data = 6'b101010;
12'b10101011000011: data = 6'b101010;
12'b10101011000100: data = 6'b101010;
12'b10101011000101: data = 6'b101010;
12'b10101011000110: data = 6'b101010;
12'b10101011000111: data = 6'b101010;
12'b10101011001000: data = 6'b101010;
12'b10101011001001: data = 6'b101010;
12'b10101011001010: data = 6'b101010;
12'b10101011001011: data = 6'b101010;
12'b10101011001100: data = 6'b101010;
12'b10101011001101: data = 6'b101010;
12'b10101011001110: data = 6'b101010;
12'b10101011001111: data = 6'b101010;
12'b10101011010000: data = 6'b101010;
12'b10101011010001: data = 6'b101010;
12'b10101011010010: data = 6'b101010;
12'b10101011010011: data = 6'b101010;
12'b10101011010100: data = 6'b101010;
12'b10101011010101: data = 6'b101010;
12'b10101011010110: data = 6'b101010;
12'b10101011010111: data = 6'b101010;
12'b10101011011000: data = 6'b101010;
12'b10101011011001: data = 6'b101010;
12'b10101011011010: data = 6'b101010;
12'b10101011011011: data = 6'b101010;
12'b10101011011100: data = 6'b101010;
12'b10101011011101: data = 6'b101010;
12'b10101011011110: data = 6'b101010;
12'b10101011011111: data = 6'b101010;
12'b10101011100000: data = 6'b101010;
12'b10101011100001: data = 6'b101010;
12'b10101011100010: data = 6'b101010;
12'b10101011100011: data = 6'b101010;
12'b10101011100100: data = 6'b101010;
12'b10101011100101: data = 6'b101010;
12'b10101011100110: data = 6'b101010;
12'b10101011100111: data = 6'b101010;
12'b10101011101000: data = 6'b101010;
12'b10101011101001: data = 6'b101010;
12'b10101011101010: data = 6'b101010;
12'b10101011101011: data = 6'b101010;
12'b10101011101100: data = 6'b101010;
12'b10101011101101: data = 6'b101010;
12'b10101011101110: data = 6'b101010;
12'b10101011101111: data = 6'b101010;
12'b10101011110000: data = 6'b101010;
12'b10101011110001: data = 6'b101010;
12'b10101011110010: data = 6'b101010;
12'b10101011110011: data = 6'b101010;
12'b10101011110100: data = 6'b101010;
12'b10101011110101: data = 6'b101010;
12'b10101011110110: data = 6'b101010;
12'b10101011110111: data = 6'b101010;
12'b10101011111000: data = 6'b101010;
12'b10101011111001: data = 6'b101010;
12'b10101011111010: data = 6'b101010;
12'b10101011111011: data = 6'b101010;
12'b10101011111100: data = 6'b101010;
12'b10101011111101: data = 6'b101010;
12'b10101011111110: data = 6'b101010;
12'b10101011111111: data = 6'b101010;
12'b101010110000000: data = 6'b101010;
12'b101010110000001: data = 6'b101010;
12'b101010110000010: data = 6'b101010;
12'b101010110000011: data = 6'b101010;
12'b101010110000100: data = 6'b101010;
12'b101010110000101: data = 6'b101010;
12'b101010110000110: data = 6'b101010;
12'b101010110000111: data = 6'b101010;
12'b101010110001000: data = 6'b101010;
12'b101010110001001: data = 6'b010101;
12'b101010110001010: data = 6'b010101;
12'b101010110001011: data = 6'b010101;
12'b101010110001100: data = 6'b000000;
12'b101010110001101: data = 6'b000000;
12'b101010110001110: data = 6'b101010;
12'b101010110001111: data = 6'b101010;
12'b101010110010000: data = 6'b101010;
12'b101010110010001: data = 6'b101010;
12'b101010110010010: data = 6'b010101;
12'b101010110010011: data = 6'b010101;
12'b101010110010100: data = 6'b010101;
12'b101010110010101: data = 6'b010101;
12'b101010110010110: data = 6'b010101;
12'b101010110010111: data = 6'b010101;
12'b101010110011000: data = 6'b010101;
12'b101010110011001: data = 6'b010101;
12'b101010110011010: data = 6'b010101;
12'b101010110011011: data = 6'b010101;
12'b101010110011100: data = 6'b010101;
12'b101010110011101: data = 6'b010101;
12'b101010110011110: data = 6'b010101;
12'b101010110011111: data = 6'b010101;
12'b101010110100000: data = 6'b010101;
12'b101010110100001: data = 6'b010101;
12'b101010110100010: data = 6'b010101;
12'b101010110100011: data = 6'b010101;
12'b101010110100100: data = 6'b010101;
12'b101010110100101: data = 6'b010101;
12'b101010110100110: data = 6'b010101;
12'b101010110100111: data = 6'b010101;
12'b101010110101000: data = 6'b010101;
12'b101010110101001: data = 6'b010101;
12'b101010110101010: data = 6'b010101;
12'b1010110000000: data = 6'b010101;
12'b1010110000001: data = 6'b010101;
12'b1010110000010: data = 6'b010101;
12'b1010110000011: data = 6'b010101;
12'b1010110000100: data = 6'b010101;
12'b1010110000101: data = 6'b010101;
12'b1010110000110: data = 6'b010101;
12'b1010110000111: data = 6'b010101;
12'b1010110001000: data = 6'b010101;
12'b1010110001001: data = 6'b010101;
12'b1010110001010: data = 6'b010101;
12'b1010110001011: data = 6'b010101;
12'b1010110001100: data = 6'b010101;
12'b1010110001101: data = 6'b010101;
12'b1010110001110: data = 6'b010101;
12'b1010110001111: data = 6'b010101;
12'b1010110010000: data = 6'b010101;
12'b1010110010001: data = 6'b010101;
12'b1010110010010: data = 6'b010101;
12'b1010110010011: data = 6'b010101;
12'b1010110010100: data = 6'b010101;
12'b1010110010101: data = 6'b010101;
12'b1010110010110: data = 6'b010101;
12'b1010110010111: data = 6'b010101;
12'b1010110011000: data = 6'b010101;
12'b1010110011001: data = 6'b101010;
12'b1010110011010: data = 6'b101010;
12'b1010110011011: data = 6'b101010;
12'b1010110011100: data = 6'b010101;
12'b1010110011101: data = 6'b000000;
12'b1010110011110: data = 6'b000000;
12'b1010110011111: data = 6'b010101;
12'b1010110100000: data = 6'b010101;
12'b1010110100001: data = 6'b010101;
12'b1010110100010: data = 6'b101010;
12'b1010110100011: data = 6'b101010;
12'b1010110100100: data = 6'b101010;
12'b1010110100101: data = 6'b101010;
12'b1010110100110: data = 6'b101010;
12'b1010110100111: data = 6'b101010;
12'b1010110101000: data = 6'b101010;
12'b1010110101001: data = 6'b101010;
12'b1010110101010: data = 6'b101010;
12'b1010110101011: data = 6'b101010;
12'b1010110101100: data = 6'b101010;
12'b1010110101101: data = 6'b101010;
12'b1010110101110: data = 6'b101010;
12'b1010110101111: data = 6'b101010;
12'b1010110110000: data = 6'b101010;
12'b1010110110001: data = 6'b101010;
12'b1010110110010: data = 6'b101010;
12'b1010110110011: data = 6'b101010;
12'b1010110110100: data = 6'b101010;
12'b1010110110101: data = 6'b101010;
12'b1010110110110: data = 6'b101010;
12'b1010110110111: data = 6'b101010;
12'b1010110111000: data = 6'b101010;
12'b1010110111001: data = 6'b101010;
12'b1010110111010: data = 6'b101010;
12'b1010110111011: data = 6'b101010;
12'b1010110111100: data = 6'b101010;
12'b1010110111101: data = 6'b101010;
12'b1010110111110: data = 6'b101010;
12'b1010110111111: data = 6'b101010;
12'b10101101000000: data = 6'b101010;
12'b10101101000001: data = 6'b101010;
12'b10101101000010: data = 6'b101010;
12'b10101101000011: data = 6'b101010;
12'b10101101000100: data = 6'b101010;
12'b10101101000101: data = 6'b101010;
12'b10101101000110: data = 6'b101010;
12'b10101101000111: data = 6'b101010;
12'b10101101001000: data = 6'b101010;
12'b10101101001001: data = 6'b101010;
12'b10101101001010: data = 6'b101010;
12'b10101101001011: data = 6'b101010;
12'b10101101001100: data = 6'b101010;
12'b10101101001101: data = 6'b101010;
12'b10101101001110: data = 6'b101010;
12'b10101101001111: data = 6'b101010;
12'b10101101010000: data = 6'b101010;
12'b10101101010001: data = 6'b101010;
12'b10101101010010: data = 6'b101010;
12'b10101101010011: data = 6'b101010;
12'b10101101010100: data = 6'b101010;
12'b10101101010101: data = 6'b101010;
12'b10101101010110: data = 6'b101010;
12'b10101101010111: data = 6'b101010;
12'b10101101011000: data = 6'b101010;
12'b10101101011001: data = 6'b101010;
12'b10101101011010: data = 6'b101010;
12'b10101101011011: data = 6'b101010;
12'b10101101011100: data = 6'b101010;
12'b10101101011101: data = 6'b101010;
12'b10101101011110: data = 6'b101010;
12'b10101101011111: data = 6'b101010;
12'b10101101100000: data = 6'b101010;
12'b10101101100001: data = 6'b101010;
12'b10101101100010: data = 6'b101010;
12'b10101101100011: data = 6'b101010;
12'b10101101100100: data = 6'b101010;
12'b10101101100101: data = 6'b101010;
12'b10101101100110: data = 6'b101010;
12'b10101101100111: data = 6'b101010;
12'b10101101101000: data = 6'b101010;
12'b10101101101001: data = 6'b101010;
12'b10101101101010: data = 6'b101010;
12'b10101101101011: data = 6'b101010;
12'b10101101101100: data = 6'b101010;
12'b10101101101101: data = 6'b101010;
12'b10101101101110: data = 6'b101010;
12'b10101101101111: data = 6'b101010;
12'b10101101110000: data = 6'b101010;
12'b10101101110001: data = 6'b101010;
12'b10101101110010: data = 6'b101010;
12'b10101101110011: data = 6'b101010;
12'b10101101110100: data = 6'b101010;
12'b10101101110101: data = 6'b101010;
12'b10101101110110: data = 6'b101010;
12'b10101101110111: data = 6'b101010;
12'b10101101111000: data = 6'b101010;
12'b10101101111001: data = 6'b101010;
12'b10101101111010: data = 6'b101010;
12'b10101101111011: data = 6'b101010;
12'b10101101111100: data = 6'b101010;
12'b10101101111101: data = 6'b101010;
12'b10101101111110: data = 6'b101010;
12'b10101101111111: data = 6'b101010;
12'b101011010000000: data = 6'b101010;
12'b101011010000001: data = 6'b101010;
12'b101011010000010: data = 6'b101010;
12'b101011010000011: data = 6'b101010;
12'b101011010000100: data = 6'b101010;
12'b101011010000101: data = 6'b101010;
12'b101011010000110: data = 6'b101010;
12'b101011010000111: data = 6'b101010;
12'b101011010001000: data = 6'b101010;
12'b101011010001001: data = 6'b010101;
12'b101011010001010: data = 6'b010101;
12'b101011010001011: data = 6'b010101;
12'b101011010001100: data = 6'b000000;
12'b101011010001101: data = 6'b000000;
12'b101011010001110: data = 6'b101010;
12'b101011010001111: data = 6'b101010;
12'b101011010010000: data = 6'b101010;
12'b101011010010001: data = 6'b101010;
12'b101011010010010: data = 6'b010101;
12'b101011010010011: data = 6'b010101;
12'b101011010010100: data = 6'b010101;
12'b101011010010101: data = 6'b010101;
12'b101011010010110: data = 6'b010101;
12'b101011010010111: data = 6'b010101;
12'b101011010011000: data = 6'b010101;
12'b101011010011001: data = 6'b010101;
12'b101011010011010: data = 6'b010101;
12'b101011010011011: data = 6'b010101;
12'b101011010011100: data = 6'b010101;
12'b101011010011101: data = 6'b010101;
12'b101011010011110: data = 6'b010101;
12'b101011010011111: data = 6'b010101;
12'b101011010100000: data = 6'b010101;
12'b101011010100001: data = 6'b010101;
12'b101011010100010: data = 6'b010101;
12'b101011010100011: data = 6'b010101;
12'b101011010100100: data = 6'b010101;
12'b101011010100101: data = 6'b010101;
12'b101011010100110: data = 6'b010101;
12'b101011010100111: data = 6'b010101;
12'b101011010101000: data = 6'b010101;
12'b101011010101001: data = 6'b010101;
12'b101011010101010: data = 6'b010101;
12'b1010111000000: data = 6'b010101;
12'b1010111000001: data = 6'b010101;
12'b1010111000010: data = 6'b010101;
12'b1010111000011: data = 6'b010101;
12'b1010111000100: data = 6'b010101;
12'b1010111000101: data = 6'b010101;
12'b1010111000110: data = 6'b010101;
12'b1010111000111: data = 6'b010101;
12'b1010111001000: data = 6'b010101;
12'b1010111001001: data = 6'b010101;
12'b1010111001010: data = 6'b010101;
12'b1010111001011: data = 6'b010101;
12'b1010111001100: data = 6'b010101;
12'b1010111001101: data = 6'b010101;
12'b1010111001110: data = 6'b010101;
12'b1010111001111: data = 6'b010101;
12'b1010111010000: data = 6'b010101;
12'b1010111010001: data = 6'b010101;
12'b1010111010010: data = 6'b010101;
12'b1010111010011: data = 6'b010101;
12'b1010111010100: data = 6'b010101;
12'b1010111010101: data = 6'b010101;
12'b1010111010110: data = 6'b010101;
12'b1010111010111: data = 6'b010101;
12'b1010111011000: data = 6'b010101;
12'b1010111011001: data = 6'b101010;
12'b1010111011010: data = 6'b101010;
12'b1010111011011: data = 6'b101010;
12'b1010111011100: data = 6'b010101;
12'b1010111011101: data = 6'b000000;
12'b1010111011110: data = 6'b000000;
12'b1010111011111: data = 6'b010101;
12'b1010111100000: data = 6'b010101;
12'b1010111100001: data = 6'b010101;
12'b1010111100010: data = 6'b101010;
12'b1010111100011: data = 6'b101010;
12'b1010111100100: data = 6'b101010;
12'b1010111100101: data = 6'b101010;
12'b1010111100110: data = 6'b101010;
12'b1010111100111: data = 6'b101010;
12'b1010111101000: data = 6'b101010;
12'b1010111101001: data = 6'b101010;
12'b1010111101010: data = 6'b101010;
12'b1010111101011: data = 6'b101010;
12'b1010111101100: data = 6'b101010;
12'b1010111101101: data = 6'b101010;
12'b1010111101110: data = 6'b101010;
12'b1010111101111: data = 6'b101010;
12'b1010111110000: data = 6'b101010;
12'b1010111110001: data = 6'b101010;
12'b1010111110010: data = 6'b101010;
12'b1010111110011: data = 6'b101010;
12'b1010111110100: data = 6'b101010;
12'b1010111110101: data = 6'b101010;
12'b1010111110110: data = 6'b101010;
12'b1010111110111: data = 6'b101010;
12'b1010111111000: data = 6'b101010;
12'b1010111111001: data = 6'b101010;
12'b1010111111010: data = 6'b101010;
12'b1010111111011: data = 6'b101010;
12'b1010111111100: data = 6'b101010;
12'b1010111111101: data = 6'b101010;
12'b1010111111110: data = 6'b101010;
12'b1010111111111: data = 6'b101010;
12'b10101111000000: data = 6'b101010;
12'b10101111000001: data = 6'b101010;
12'b10101111000010: data = 6'b101010;
12'b10101111000011: data = 6'b101010;
12'b10101111000100: data = 6'b101010;
12'b10101111000101: data = 6'b101010;
12'b10101111000110: data = 6'b101010;
12'b10101111000111: data = 6'b101010;
12'b10101111001000: data = 6'b101010;
12'b10101111001001: data = 6'b101010;
12'b10101111001010: data = 6'b101010;
12'b10101111001011: data = 6'b101010;
12'b10101111001100: data = 6'b101010;
12'b10101111001101: data = 6'b101010;
12'b10101111001110: data = 6'b101010;
12'b10101111001111: data = 6'b101010;
12'b10101111010000: data = 6'b101010;
12'b10101111010001: data = 6'b101010;
12'b10101111010010: data = 6'b101010;
12'b10101111010011: data = 6'b101010;
12'b10101111010100: data = 6'b101010;
12'b10101111010101: data = 6'b101010;
12'b10101111010110: data = 6'b101010;
12'b10101111010111: data = 6'b101010;
12'b10101111011000: data = 6'b101010;
12'b10101111011001: data = 6'b101010;
12'b10101111011010: data = 6'b101010;
12'b10101111011011: data = 6'b101010;
12'b10101111011100: data = 6'b101010;
12'b10101111011101: data = 6'b101010;
12'b10101111011110: data = 6'b101010;
12'b10101111011111: data = 6'b101010;
12'b10101111100000: data = 6'b101010;
12'b10101111100001: data = 6'b101010;
12'b10101111100010: data = 6'b101010;
12'b10101111100011: data = 6'b101010;
12'b10101111100100: data = 6'b101010;
12'b10101111100101: data = 6'b101010;
12'b10101111100110: data = 6'b101010;
12'b10101111100111: data = 6'b101010;
12'b10101111101000: data = 6'b101010;
12'b10101111101001: data = 6'b101010;
12'b10101111101010: data = 6'b101010;
12'b10101111101011: data = 6'b101010;
12'b10101111101100: data = 6'b101010;
12'b10101111101101: data = 6'b101010;
12'b10101111101110: data = 6'b101010;
12'b10101111101111: data = 6'b101010;
12'b10101111110000: data = 6'b101010;
12'b10101111110001: data = 6'b101010;
12'b10101111110010: data = 6'b101010;
12'b10101111110011: data = 6'b101010;
12'b10101111110100: data = 6'b101010;
12'b10101111110101: data = 6'b101010;
12'b10101111110110: data = 6'b101010;
12'b10101111110111: data = 6'b101010;
12'b10101111111000: data = 6'b101010;
12'b10101111111001: data = 6'b101010;
12'b10101111111010: data = 6'b101010;
12'b10101111111011: data = 6'b101010;
12'b10101111111100: data = 6'b101010;
12'b10101111111101: data = 6'b101010;
12'b10101111111110: data = 6'b101010;
12'b10101111111111: data = 6'b101010;
12'b101011110000000: data = 6'b101010;
12'b101011110000001: data = 6'b101010;
12'b101011110000010: data = 6'b101010;
12'b101011110000011: data = 6'b101010;
12'b101011110000100: data = 6'b101010;
12'b101011110000101: data = 6'b101010;
12'b101011110000110: data = 6'b101010;
12'b101011110000111: data = 6'b101010;
12'b101011110001000: data = 6'b101010;
12'b101011110001001: data = 6'b010101;
12'b101011110001010: data = 6'b010101;
12'b101011110001011: data = 6'b010101;
12'b101011110001100: data = 6'b000000;
12'b101011110001101: data = 6'b000000;
12'b101011110001110: data = 6'b101010;
12'b101011110001111: data = 6'b101010;
12'b101011110010000: data = 6'b101010;
12'b101011110010001: data = 6'b101010;
12'b101011110010010: data = 6'b010101;
12'b101011110010011: data = 6'b010101;
12'b101011110010100: data = 6'b010101;
12'b101011110010101: data = 6'b010101;
12'b101011110010110: data = 6'b010101;
12'b101011110010111: data = 6'b010101;
12'b101011110011000: data = 6'b010101;
12'b101011110011001: data = 6'b010101;
12'b101011110011010: data = 6'b010101;
12'b101011110011011: data = 6'b010101;
12'b101011110011100: data = 6'b010101;
12'b101011110011101: data = 6'b010101;
12'b101011110011110: data = 6'b010101;
12'b101011110011111: data = 6'b010101;
12'b101011110100000: data = 6'b010101;
12'b101011110100001: data = 6'b010101;
12'b101011110100010: data = 6'b010101;
12'b101011110100011: data = 6'b010101;
12'b101011110100100: data = 6'b010101;
12'b101011110100101: data = 6'b010101;
12'b101011110100110: data = 6'b010101;
12'b101011110100111: data = 6'b010101;
12'b101011110101000: data = 6'b010101;
12'b101011110101001: data = 6'b010101;
12'b101011110101010: data = 6'b010101;
12'b1011000000000: data = 6'b010101;
12'b1011000000001: data = 6'b010101;
12'b1011000000010: data = 6'b010101;
12'b1011000000011: data = 6'b010101;
12'b1011000000100: data = 6'b010101;
12'b1011000000101: data = 6'b010101;
12'b1011000000110: data = 6'b010101;
12'b1011000000111: data = 6'b010101;
12'b1011000001000: data = 6'b010101;
12'b1011000001001: data = 6'b010101;
12'b1011000001010: data = 6'b010101;
12'b1011000001011: data = 6'b010101;
12'b1011000001100: data = 6'b010101;
12'b1011000001101: data = 6'b010101;
12'b1011000001110: data = 6'b010101;
12'b1011000001111: data = 6'b010101;
12'b1011000010000: data = 6'b010101;
12'b1011000010001: data = 6'b010101;
12'b1011000010010: data = 6'b010101;
12'b1011000010011: data = 6'b010101;
12'b1011000010100: data = 6'b010101;
12'b1011000010101: data = 6'b010101;
12'b1011000010110: data = 6'b010101;
12'b1011000010111: data = 6'b010101;
12'b1011000011000: data = 6'b010101;
12'b1011000011001: data = 6'b101010;
12'b1011000011010: data = 6'b101010;
12'b1011000011011: data = 6'b101010;
12'b1011000011100: data = 6'b010101;
12'b1011000011101: data = 6'b000000;
12'b1011000011110: data = 6'b000000;
12'b1011000011111: data = 6'b010101;
12'b1011000100000: data = 6'b010101;
12'b1011000100001: data = 6'b010101;
12'b1011000100010: data = 6'b010101;
12'b1011000100011: data = 6'b101001;
12'b1011000100100: data = 6'b101010;
12'b1011000100101: data = 6'b101010;
12'b1011000100110: data = 6'b101010;
12'b1011000100111: data = 6'b101010;
12'b1011000101000: data = 6'b101010;
12'b1011000101001: data = 6'b101010;
12'b1011000101010: data = 6'b101010;
12'b1011000101011: data = 6'b101010;
12'b1011000101100: data = 6'b101010;
12'b1011000101101: data = 6'b101010;
12'b1011000101110: data = 6'b101010;
12'b1011000101111: data = 6'b101010;
12'b1011000110000: data = 6'b101010;
12'b1011000110001: data = 6'b101010;
12'b1011000110010: data = 6'b101010;
12'b1011000110011: data = 6'b101010;
12'b1011000110100: data = 6'b101010;
12'b1011000110101: data = 6'b101010;
12'b1011000110110: data = 6'b101010;
12'b1011000110111: data = 6'b101010;
12'b1011000111000: data = 6'b101010;
12'b1011000111001: data = 6'b101010;
12'b1011000111010: data = 6'b101010;
12'b1011000111011: data = 6'b101010;
12'b1011000111100: data = 6'b111110;
12'b1011000111101: data = 6'b111110;
12'b1011000111110: data = 6'b111110;
12'b1011000111111: data = 6'b111110;
12'b10110001000000: data = 6'b111110;
12'b10110001000001: data = 6'b111110;
12'b10110001000010: data = 6'b111110;
12'b10110001000011: data = 6'b111110;
12'b10110001000100: data = 6'b111110;
12'b10110001000101: data = 6'b101010;
12'b10110001000110: data = 6'b101010;
12'b10110001000111: data = 6'b111010;
12'b10110001001000: data = 6'b111010;
12'b10110001001001: data = 6'b101010;
12'b10110001001010: data = 6'b101010;
12'b10110001001011: data = 6'b101010;
12'b10110001001100: data = 6'b101010;
12'b10110001001101: data = 6'b101010;
12'b10110001001110: data = 6'b101010;
12'b10110001001111: data = 6'b101010;
12'b10110001010000: data = 6'b101010;
12'b10110001010001: data = 6'b101010;
12'b10110001010010: data = 6'b101010;
12'b10110001010011: data = 6'b101010;
12'b10110001010100: data = 6'b101010;
12'b10110001010101: data = 6'b101010;
12'b10110001010110: data = 6'b101010;
12'b10110001010111: data = 6'b101010;
12'b10110001011000: data = 6'b101010;
12'b10110001011001: data = 6'b101010;
12'b10110001011010: data = 6'b101010;
12'b10110001011011: data = 6'b101010;
12'b10110001011100: data = 6'b101010;
12'b10110001011101: data = 6'b101010;
12'b10110001011110: data = 6'b101010;
12'b10110001011111: data = 6'b101010;
12'b10110001100000: data = 6'b101010;
12'b10110001100001: data = 6'b101010;
12'b10110001100010: data = 6'b101010;
12'b10110001100011: data = 6'b101010;
12'b10110001100100: data = 6'b101010;
12'b10110001100101: data = 6'b101010;
12'b10110001100110: data = 6'b101010;
12'b10110001100111: data = 6'b101010;
12'b10110001101000: data = 6'b101010;
12'b10110001101001: data = 6'b101010;
12'b10110001101010: data = 6'b101010;
12'b10110001101011: data = 6'b101010;
12'b10110001101100: data = 6'b101010;
12'b10110001101101: data = 6'b101010;
12'b10110001101110: data = 6'b101010;
12'b10110001101111: data = 6'b101010;
12'b10110001110000: data = 6'b101010;
12'b10110001110001: data = 6'b101010;
12'b10110001110010: data = 6'b101010;
12'b10110001110011: data = 6'b101010;
12'b10110001110100: data = 6'b101010;
12'b10110001110101: data = 6'b101010;
12'b10110001110110: data = 6'b101010;
12'b10110001110111: data = 6'b101010;
12'b10110001111000: data = 6'b101010;
12'b10110001111001: data = 6'b101010;
12'b10110001111010: data = 6'b101010;
12'b10110001111011: data = 6'b101010;
12'b10110001111100: data = 6'b101010;
12'b10110001111101: data = 6'b101010;
12'b10110001111110: data = 6'b101010;
12'b10110001111111: data = 6'b101010;
12'b101100010000000: data = 6'b101010;
12'b101100010000001: data = 6'b101010;
12'b101100010000010: data = 6'b101010;
12'b101100010000011: data = 6'b101010;
12'b101100010000100: data = 6'b101010;
12'b101100010000101: data = 6'b101010;
12'b101100010000110: data = 6'b010101;
12'b101100010000111: data = 6'b010101;
12'b101100010001000: data = 6'b010101;
12'b101100010001001: data = 6'b010101;
12'b101100010001010: data = 6'b010101;
12'b101100010001011: data = 6'b010101;
12'b101100010001100: data = 6'b000000;
12'b101100010001101: data = 6'b000000;
12'b101100010001110: data = 6'b101010;
12'b101100010001111: data = 6'b101010;
12'b101100010010000: data = 6'b101010;
12'b101100010010001: data = 6'b101010;
12'b101100010010010: data = 6'b010101;
12'b101100010010011: data = 6'b010101;
12'b101100010010100: data = 6'b010101;
12'b101100010010101: data = 6'b010101;
12'b101100010010110: data = 6'b010101;
12'b101100010010111: data = 6'b010101;
12'b101100010011000: data = 6'b010101;
12'b101100010011001: data = 6'b010101;
12'b101100010011010: data = 6'b010101;
12'b101100010011011: data = 6'b010101;
12'b101100010011100: data = 6'b010101;
12'b101100010011101: data = 6'b010101;
12'b101100010011110: data = 6'b010101;
12'b101100010011111: data = 6'b010101;
12'b101100010100000: data = 6'b010101;
12'b101100010100001: data = 6'b010101;
12'b101100010100010: data = 6'b010101;
12'b101100010100011: data = 6'b010101;
12'b101100010100100: data = 6'b010101;
12'b101100010100101: data = 6'b010101;
12'b101100010100110: data = 6'b010101;
12'b101100010100111: data = 6'b010101;
12'b101100010101000: data = 6'b010101;
12'b101100010101001: data = 6'b010101;
12'b101100010101010: data = 6'b010101;
12'b1011001000000: data = 6'b010101;
12'b1011001000001: data = 6'b010101;
12'b1011001000010: data = 6'b010101;
12'b1011001000011: data = 6'b010101;
12'b1011001000100: data = 6'b010101;
12'b1011001000101: data = 6'b010101;
12'b1011001000110: data = 6'b010101;
12'b1011001000111: data = 6'b010101;
12'b1011001001000: data = 6'b010101;
12'b1011001001001: data = 6'b010101;
12'b1011001001010: data = 6'b010101;
12'b1011001001011: data = 6'b010101;
12'b1011001001100: data = 6'b010101;
12'b1011001001101: data = 6'b010101;
12'b1011001001110: data = 6'b010101;
12'b1011001001111: data = 6'b010101;
12'b1011001010000: data = 6'b010101;
12'b1011001010001: data = 6'b010101;
12'b1011001010010: data = 6'b010101;
12'b1011001010011: data = 6'b010101;
12'b1011001010100: data = 6'b010101;
12'b1011001010101: data = 6'b010101;
12'b1011001010110: data = 6'b010101;
12'b1011001010111: data = 6'b010101;
12'b1011001011000: data = 6'b010101;
12'b1011001011001: data = 6'b101010;
12'b1011001011010: data = 6'b101010;
12'b1011001011011: data = 6'b101010;
12'b1011001011100: data = 6'b010101;
12'b1011001011101: data = 6'b000000;
12'b1011001011110: data = 6'b000000;
12'b1011001011111: data = 6'b010101;
12'b1011001100000: data = 6'b010101;
12'b1011001100001: data = 6'b010101;
12'b1011001100010: data = 6'b010101;
12'b1011001100011: data = 6'b010101;
12'b1011001100100: data = 6'b010101;
12'b1011001100101: data = 6'b101010;
12'b1011001100110: data = 6'b101010;
12'b1011001100111: data = 6'b101010;
12'b1011001101000: data = 6'b101010;
12'b1011001101001: data = 6'b101010;
12'b1011001101010: data = 6'b101010;
12'b1011001101011: data = 6'b101010;
12'b1011001101100: data = 6'b101010;
12'b1011001101101: data = 6'b101010;
12'b1011001101110: data = 6'b101010;
12'b1011001101111: data = 6'b101010;
12'b1011001110000: data = 6'b101010;
12'b1011001110001: data = 6'b101010;
12'b1011001110010: data = 6'b101010;
12'b1011001110011: data = 6'b101010;
12'b1011001110100: data = 6'b101010;
12'b1011001110101: data = 6'b101010;
12'b1011001110110: data = 6'b101010;
12'b1011001110111: data = 6'b101010;
12'b1011001111000: data = 6'b111110;
12'b1011001111001: data = 6'b111110;
12'b1011001111010: data = 6'b111110;
12'b1011001111011: data = 6'b111110;
12'b1011001111100: data = 6'b111111;
12'b1011001111101: data = 6'b111111;
12'b1011001111110: data = 6'b111111;
12'b1011001111111: data = 6'b111111;
12'b10110011000000: data = 6'b111111;
12'b10110011000001: data = 6'b111111;
12'b10110011000010: data = 6'b111111;
12'b10110011000011: data = 6'b111110;
12'b10110011000100: data = 6'b111110;
12'b10110011000101: data = 6'b111110;
12'b10110011000110: data = 6'b111110;
12'b10110011000111: data = 6'b111110;
12'b10110011001000: data = 6'b111110;
12'b10110011001001: data = 6'b111110;
12'b10110011001010: data = 6'b101010;
12'b10110011001011: data = 6'b111110;
12'b10110011001100: data = 6'b111010;
12'b10110011001101: data = 6'b101010;
12'b10110011001110: data = 6'b111010;
12'b10110011001111: data = 6'b101010;
12'b10110011010000: data = 6'b101010;
12'b10110011010001: data = 6'b101010;
12'b10110011010010: data = 6'b101010;
12'b10110011010011: data = 6'b101010;
12'b10110011010100: data = 6'b101010;
12'b10110011010101: data = 6'b101010;
12'b10110011010110: data = 6'b101010;
12'b10110011010111: data = 6'b101010;
12'b10110011011000: data = 6'b101010;
12'b10110011011001: data = 6'b101010;
12'b10110011011010: data = 6'b101010;
12'b10110011011011: data = 6'b101010;
12'b10110011011100: data = 6'b101010;
12'b10110011011101: data = 6'b101010;
12'b10110011011110: data = 6'b101010;
12'b10110011011111: data = 6'b101010;
12'b10110011100000: data = 6'b101010;
12'b10110011100001: data = 6'b101010;
12'b10110011100010: data = 6'b101010;
12'b10110011100011: data = 6'b101010;
12'b10110011100100: data = 6'b101010;
12'b10110011100101: data = 6'b101010;
12'b10110011100110: data = 6'b101010;
12'b10110011100111: data = 6'b101010;
12'b10110011101000: data = 6'b101010;
12'b10110011101001: data = 6'b101010;
12'b10110011101010: data = 6'b101010;
12'b10110011101011: data = 6'b101010;
12'b10110011101100: data = 6'b101010;
12'b10110011101101: data = 6'b101010;
12'b10110011101110: data = 6'b101010;
12'b10110011101111: data = 6'b101010;
12'b10110011110000: data = 6'b101010;
12'b10110011110001: data = 6'b101010;
12'b10110011110010: data = 6'b101010;
12'b10110011110011: data = 6'b101010;
12'b10110011110100: data = 6'b101010;
12'b10110011110101: data = 6'b101010;
12'b10110011110110: data = 6'b101010;
12'b10110011110111: data = 6'b101010;
12'b10110011111000: data = 6'b101010;
12'b10110011111001: data = 6'b101010;
12'b10110011111010: data = 6'b101010;
12'b10110011111011: data = 6'b101010;
12'b10110011111100: data = 6'b101010;
12'b10110011111101: data = 6'b101010;
12'b10110011111110: data = 6'b101010;
12'b10110011111111: data = 6'b101010;
12'b101100110000000: data = 6'b101010;
12'b101100110000001: data = 6'b101010;
12'b101100110000010: data = 6'b101010;
12'b101100110000011: data = 6'b101010;
12'b101100110000100: data = 6'b101010;
12'b101100110000101: data = 6'b101010;
12'b101100110000110: data = 6'b010101;
12'b101100110000111: data = 6'b010101;
12'b101100110001000: data = 6'b010101;
12'b101100110001001: data = 6'b010101;
12'b101100110001010: data = 6'b010101;
12'b101100110001011: data = 6'b010101;
12'b101100110001100: data = 6'b000000;
12'b101100110001101: data = 6'b000000;
12'b101100110001110: data = 6'b101010;
12'b101100110001111: data = 6'b101010;
12'b101100110010000: data = 6'b101010;
12'b101100110010001: data = 6'b101010;
12'b101100110010010: data = 6'b010101;
12'b101100110010011: data = 6'b010101;
12'b101100110010100: data = 6'b010101;
12'b101100110010101: data = 6'b010101;
12'b101100110010110: data = 6'b010101;
12'b101100110010111: data = 6'b010101;
12'b101100110011000: data = 6'b010101;
12'b101100110011001: data = 6'b010101;
12'b101100110011010: data = 6'b010101;
12'b101100110011011: data = 6'b010101;
12'b101100110011100: data = 6'b010101;
12'b101100110011101: data = 6'b010101;
12'b101100110011110: data = 6'b010101;
12'b101100110011111: data = 6'b010101;
12'b101100110100000: data = 6'b010101;
12'b101100110100001: data = 6'b010101;
12'b101100110100010: data = 6'b010101;
12'b101100110100011: data = 6'b010101;
12'b101100110100100: data = 6'b010101;
12'b101100110100101: data = 6'b010101;
12'b101100110100110: data = 6'b010101;
12'b101100110100111: data = 6'b010101;
12'b101100110101000: data = 6'b010101;
12'b101100110101001: data = 6'b010101;
12'b101100110101010: data = 6'b010101;
12'b1011010000000: data = 6'b010101;
12'b1011010000001: data = 6'b010101;
12'b1011010000010: data = 6'b010101;
12'b1011010000011: data = 6'b010101;
12'b1011010000100: data = 6'b010101;
12'b1011010000101: data = 6'b010101;
12'b1011010000110: data = 6'b010101;
12'b1011010000111: data = 6'b010101;
12'b1011010001000: data = 6'b010101;
12'b1011010001001: data = 6'b010101;
12'b1011010001010: data = 6'b010101;
12'b1011010001011: data = 6'b010101;
12'b1011010001100: data = 6'b010101;
12'b1011010001101: data = 6'b010101;
12'b1011010001110: data = 6'b010101;
12'b1011010001111: data = 6'b010101;
12'b1011010010000: data = 6'b010101;
12'b1011010010001: data = 6'b010101;
12'b1011010010010: data = 6'b010101;
12'b1011010010011: data = 6'b010101;
12'b1011010010100: data = 6'b010101;
12'b1011010010101: data = 6'b010101;
12'b1011010010110: data = 6'b010101;
12'b1011010010111: data = 6'b010101;
12'b1011010011000: data = 6'b010101;
12'b1011010011001: data = 6'b101010;
12'b1011010011010: data = 6'b101010;
12'b1011010011011: data = 6'b101010;
12'b1011010011100: data = 6'b010101;
12'b1011010011101: data = 6'b000000;
12'b1011010011110: data = 6'b000000;
12'b1011010011111: data = 6'b010101;
12'b1011010100000: data = 6'b010101;
12'b1011010100001: data = 6'b010101;
12'b1011010100010: data = 6'b010101;
12'b1011010100011: data = 6'b010101;
12'b1011010100100: data = 6'b010101;
12'b1011010100101: data = 6'b101010;
12'b1011010100110: data = 6'b101010;
12'b1011010100111: data = 6'b101010;
12'b1011010101000: data = 6'b101010;
12'b1011010101001: data = 6'b101010;
12'b1011010101010: data = 6'b101010;
12'b1011010101011: data = 6'b101010;
12'b1011010101100: data = 6'b101010;
12'b1011010101101: data = 6'b101010;
12'b1011010101110: data = 6'b101010;
12'b1011010101111: data = 6'b101010;
12'b1011010110000: data = 6'b101010;
12'b1011010110001: data = 6'b101010;
12'b1011010110010: data = 6'b101010;
12'b1011010110011: data = 6'b101010;
12'b1011010110100: data = 6'b101010;
12'b1011010110101: data = 6'b101010;
12'b1011010110110: data = 6'b111010;
12'b1011010110111: data = 6'b111110;
12'b1011010111000: data = 6'b111110;
12'b1011010111001: data = 6'b111110;
12'b1011010111010: data = 6'b111111;
12'b1011010111011: data = 6'b111111;
12'b1011010111100: data = 6'b111111;
12'b1011010111101: data = 6'b111111;
12'b1011010111110: data = 6'b111111;
12'b1011010111111: data = 6'b111111;
12'b10110101000000: data = 6'b111111;
12'b10110101000001: data = 6'b111111;
12'b10110101000010: data = 6'b111111;
12'b10110101000011: data = 6'b111111;
12'b10110101000100: data = 6'b111111;
12'b10110101000101: data = 6'b111110;
12'b10110101000110: data = 6'b111110;
12'b10110101000111: data = 6'b111110;
12'b10110101001000: data = 6'b111110;
12'b10110101001001: data = 6'b111110;
12'b10110101001010: data = 6'b111010;
12'b10110101001011: data = 6'b111110;
12'b10110101001100: data = 6'b111010;
12'b10110101001101: data = 6'b111010;
12'b10110101001110: data = 6'b111010;
12'b10110101001111: data = 6'b101010;
12'b10110101010000: data = 6'b101010;
12'b10110101010001: data = 6'b101010;
12'b10110101010010: data = 6'b101010;
12'b10110101010011: data = 6'b101010;
12'b10110101010100: data = 6'b101010;
12'b10110101010101: data = 6'b101010;
12'b10110101010110: data = 6'b101010;
12'b10110101010111: data = 6'b101010;
12'b10110101011000: data = 6'b101010;
12'b10110101011001: data = 6'b101010;
12'b10110101011010: data = 6'b101010;
12'b10110101011011: data = 6'b101010;
12'b10110101011100: data = 6'b101010;
12'b10110101011101: data = 6'b101010;
12'b10110101011110: data = 6'b101010;
12'b10110101011111: data = 6'b101010;
12'b10110101100000: data = 6'b101010;
12'b10110101100001: data = 6'b101010;
12'b10110101100010: data = 6'b101010;
12'b10110101100011: data = 6'b101010;
12'b10110101100100: data = 6'b101010;
12'b10110101100101: data = 6'b101010;
12'b10110101100110: data = 6'b101010;
12'b10110101100111: data = 6'b101010;
12'b10110101101000: data = 6'b101010;
12'b10110101101001: data = 6'b101010;
12'b10110101101010: data = 6'b101010;
12'b10110101101011: data = 6'b101010;
12'b10110101101100: data = 6'b101010;
12'b10110101101101: data = 6'b101010;
12'b10110101101110: data = 6'b101010;
12'b10110101101111: data = 6'b101010;
12'b10110101110000: data = 6'b101010;
12'b10110101110001: data = 6'b101010;
12'b10110101110010: data = 6'b101010;
12'b10110101110011: data = 6'b101010;
12'b10110101110100: data = 6'b101010;
12'b10110101110101: data = 6'b101010;
12'b10110101110110: data = 6'b101010;
12'b10110101110111: data = 6'b101010;
12'b10110101111000: data = 6'b101010;
12'b10110101111001: data = 6'b101010;
12'b10110101111010: data = 6'b101010;
12'b10110101111011: data = 6'b101010;
12'b10110101111100: data = 6'b101010;
12'b10110101111101: data = 6'b101010;
12'b10110101111110: data = 6'b101010;
12'b10110101111111: data = 6'b101010;
12'b101101010000000: data = 6'b101001;
12'b101101010000001: data = 6'b101001;
12'b101101010000010: data = 6'b101001;
12'b101101010000011: data = 6'b010101;
12'b101101010000100: data = 6'b010101;
12'b101101010000101: data = 6'b010101;
12'b101101010000110: data = 6'b010101;
12'b101101010000111: data = 6'b010101;
12'b101101010001000: data = 6'b010101;
12'b101101010001001: data = 6'b010101;
12'b101101010001010: data = 6'b010101;
12'b101101010001011: data = 6'b010101;
12'b101101010001100: data = 6'b000000;
12'b101101010001101: data = 6'b000000;
12'b101101010001110: data = 6'b101010;
12'b101101010001111: data = 6'b101010;
12'b101101010010000: data = 6'b101010;
12'b101101010010001: data = 6'b101010;
12'b101101010010010: data = 6'b010101;
12'b101101010010011: data = 6'b010101;
12'b101101010010100: data = 6'b010101;
12'b101101010010101: data = 6'b010101;
12'b101101010010110: data = 6'b010101;
12'b101101010010111: data = 6'b010101;
12'b101101010011000: data = 6'b010101;
12'b101101010011001: data = 6'b010101;
12'b101101010011010: data = 6'b010101;
12'b101101010011011: data = 6'b010101;
12'b101101010011100: data = 6'b010101;
12'b101101010011101: data = 6'b010101;
12'b101101010011110: data = 6'b010101;
12'b101101010011111: data = 6'b010101;
12'b101101010100000: data = 6'b010101;
12'b101101010100001: data = 6'b010101;
12'b101101010100010: data = 6'b010101;
12'b101101010100011: data = 6'b010101;
12'b101101010100100: data = 6'b010101;
12'b101101010100101: data = 6'b010101;
12'b101101010100110: data = 6'b010101;
12'b101101010100111: data = 6'b010101;
12'b101101010101000: data = 6'b010101;
12'b101101010101001: data = 6'b010101;
12'b101101010101010: data = 6'b010101;
12'b1011011000000: data = 6'b010101;
12'b1011011000001: data = 6'b010101;
12'b1011011000010: data = 6'b010101;
12'b1011011000011: data = 6'b010101;
12'b1011011000100: data = 6'b010101;
12'b1011011000101: data = 6'b010101;
12'b1011011000110: data = 6'b010101;
12'b1011011000111: data = 6'b010101;
12'b1011011001000: data = 6'b010101;
12'b1011011001001: data = 6'b010101;
12'b1011011001010: data = 6'b010101;
12'b1011011001011: data = 6'b010101;
12'b1011011001100: data = 6'b010101;
12'b1011011001101: data = 6'b010101;
12'b1011011001110: data = 6'b010101;
12'b1011011001111: data = 6'b010101;
12'b1011011010000: data = 6'b010101;
12'b1011011010001: data = 6'b010101;
12'b1011011010010: data = 6'b010101;
12'b1011011010011: data = 6'b010101;
12'b1011011010100: data = 6'b010101;
12'b1011011010101: data = 6'b010101;
12'b1011011010110: data = 6'b010101;
12'b1011011010111: data = 6'b010101;
12'b1011011011000: data = 6'b010101;
12'b1011011011001: data = 6'b101010;
12'b1011011011010: data = 6'b101010;
12'b1011011011011: data = 6'b101010;
12'b1011011011100: data = 6'b010101;
12'b1011011011101: data = 6'b000000;
12'b1011011011110: data = 6'b000000;
12'b1011011011111: data = 6'b010101;
12'b1011011100000: data = 6'b010101;
12'b1011011100001: data = 6'b010101;
12'b1011011100010: data = 6'b010101;
12'b1011011100011: data = 6'b010101;
12'b1011011100100: data = 6'b010101;
12'b1011011100101: data = 6'b101001;
12'b1011011100110: data = 6'b101001;
12'b1011011100111: data = 6'b101010;
12'b1011011101000: data = 6'b101010;
12'b1011011101001: data = 6'b101010;
12'b1011011101010: data = 6'b101010;
12'b1011011101011: data = 6'b101010;
12'b1011011101100: data = 6'b101010;
12'b1011011101101: data = 6'b101010;
12'b1011011101110: data = 6'b101010;
12'b1011011101111: data = 6'b101010;
12'b1011011110000: data = 6'b101010;
12'b1011011110001: data = 6'b101010;
12'b1011011110010: data = 6'b101010;
12'b1011011110011: data = 6'b101010;
12'b1011011110100: data = 6'b101010;
12'b1011011110101: data = 6'b111010;
12'b1011011110110: data = 6'b111010;
12'b1011011110111: data = 6'b111110;
12'b1011011111000: data = 6'b111110;
12'b1011011111001: data = 6'b111111;
12'b1011011111010: data = 6'b111111;
12'b1011011111011: data = 6'b111111;
12'b1011011111100: data = 6'b111111;
12'b1011011111101: data = 6'b111111;
12'b1011011111110: data = 6'b111111;
12'b1011011111111: data = 6'b111111;
12'b10110111000000: data = 6'b111111;
12'b10110111000001: data = 6'b111111;
12'b10110111000010: data = 6'b111111;
12'b10110111000011: data = 6'b111111;
12'b10110111000100: data = 6'b111111;
12'b10110111000101: data = 6'b111111;
12'b10110111000110: data = 6'b111111;
12'b10110111000111: data = 6'b111110;
12'b10110111001000: data = 6'b111110;
12'b10110111001001: data = 6'b111110;
12'b10110111001010: data = 6'b111110;
12'b10110111001011: data = 6'b111110;
12'b10110111001100: data = 6'b111010;
12'b10110111001101: data = 6'b111010;
12'b10110111001110: data = 6'b111010;
12'b10110111001111: data = 6'b101010;
12'b10110111010000: data = 6'b101010;
12'b10110111010001: data = 6'b101010;
12'b10110111010010: data = 6'b101010;
12'b10110111010011: data = 6'b101010;
12'b10110111010100: data = 6'b101010;
12'b10110111010101: data = 6'b101010;
12'b10110111010110: data = 6'b101010;
12'b10110111010111: data = 6'b101010;
12'b10110111011000: data = 6'b101010;
12'b10110111011001: data = 6'b101010;
12'b10110111011010: data = 6'b101010;
12'b10110111011011: data = 6'b101010;
12'b10110111011100: data = 6'b101010;
12'b10110111011101: data = 6'b101010;
12'b10110111011110: data = 6'b101010;
12'b10110111011111: data = 6'b101010;
12'b10110111100000: data = 6'b101010;
12'b10110111100001: data = 6'b101010;
12'b10110111100010: data = 6'b101010;
12'b10110111100011: data = 6'b101010;
12'b10110111100100: data = 6'b101010;
12'b10110111100101: data = 6'b101010;
12'b10110111100110: data = 6'b101010;
12'b10110111100111: data = 6'b101010;
12'b10110111101000: data = 6'b101010;
12'b10110111101001: data = 6'b101010;
12'b10110111101010: data = 6'b101010;
12'b10110111101011: data = 6'b101010;
12'b10110111101100: data = 6'b101010;
12'b10110111101101: data = 6'b101010;
12'b10110111101110: data = 6'b101010;
12'b10110111101111: data = 6'b101010;
12'b10110111110000: data = 6'b101010;
12'b10110111110001: data = 6'b101010;
12'b10110111110010: data = 6'b101010;
12'b10110111110011: data = 6'b101010;
12'b10110111110100: data = 6'b101010;
12'b10110111110101: data = 6'b101010;
12'b10110111110110: data = 6'b101010;
12'b10110111110111: data = 6'b101010;
12'b10110111111000: data = 6'b101010;
12'b10110111111001: data = 6'b101001;
12'b10110111111010: data = 6'b101001;
12'b10110111111011: data = 6'b101001;
12'b10110111111100: data = 6'b010101;
12'b10110111111101: data = 6'b010101;
12'b10110111111110: data = 6'b010101;
12'b10110111111111: data = 6'b010101;
12'b101101110000000: data = 6'b010101;
12'b101101110000001: data = 6'b010101;
12'b101101110000010: data = 6'b010101;
12'b101101110000011: data = 6'b010101;
12'b101101110000100: data = 6'b010101;
12'b101101110000101: data = 6'b010101;
12'b101101110000110: data = 6'b010101;
12'b101101110000111: data = 6'b010101;
12'b101101110001000: data = 6'b010101;
12'b101101110001001: data = 6'b010101;
12'b101101110001010: data = 6'b010101;
12'b101101110001011: data = 6'b010101;
12'b101101110001100: data = 6'b000000;
12'b101101110001101: data = 6'b000000;
12'b101101110001110: data = 6'b101010;
12'b101101110001111: data = 6'b101010;
12'b101101110010000: data = 6'b101010;
12'b101101110010001: data = 6'b101010;
12'b101101110010010: data = 6'b010101;
12'b101101110010011: data = 6'b010101;
12'b101101110010100: data = 6'b010101;
12'b101101110010101: data = 6'b010101;
12'b101101110010110: data = 6'b010101;
12'b101101110010111: data = 6'b010101;
12'b101101110011000: data = 6'b010101;
12'b101101110011001: data = 6'b010101;
12'b101101110011010: data = 6'b010101;
12'b101101110011011: data = 6'b010101;
12'b101101110011100: data = 6'b010101;
12'b101101110011101: data = 6'b010101;
12'b101101110011110: data = 6'b010101;
12'b101101110011111: data = 6'b010101;
12'b101101110100000: data = 6'b010101;
12'b101101110100001: data = 6'b010101;
12'b101101110100010: data = 6'b010101;
12'b101101110100011: data = 6'b010101;
12'b101101110100100: data = 6'b010101;
12'b101101110100101: data = 6'b010101;
12'b101101110100110: data = 6'b010101;
12'b101101110100111: data = 6'b010101;
12'b101101110101000: data = 6'b010101;
12'b101101110101001: data = 6'b010101;
12'b101101110101010: data = 6'b010101;
12'b1011100000000: data = 6'b010101;
12'b1011100000001: data = 6'b010101;
12'b1011100000010: data = 6'b010101;
12'b1011100000011: data = 6'b010101;
12'b1011100000100: data = 6'b010101;
12'b1011100000101: data = 6'b010101;
12'b1011100000110: data = 6'b010101;
12'b1011100000111: data = 6'b010101;
12'b1011100001000: data = 6'b010101;
12'b1011100001001: data = 6'b010101;
12'b1011100001010: data = 6'b010101;
12'b1011100001011: data = 6'b010101;
12'b1011100001100: data = 6'b010101;
12'b1011100001101: data = 6'b010101;
12'b1011100001110: data = 6'b010101;
12'b1011100001111: data = 6'b010101;
12'b1011100010000: data = 6'b010101;
12'b1011100010001: data = 6'b010101;
12'b1011100010010: data = 6'b010101;
12'b1011100010011: data = 6'b010101;
12'b1011100010100: data = 6'b010101;
12'b1011100010101: data = 6'b010101;
12'b1011100010110: data = 6'b010101;
12'b1011100010111: data = 6'b010101;
12'b1011100011000: data = 6'b010101;
12'b1011100011001: data = 6'b101010;
12'b1011100011010: data = 6'b101010;
12'b1011100011011: data = 6'b101010;
12'b1011100011100: data = 6'b010101;
12'b1011100011101: data = 6'b000000;
12'b1011100011110: data = 6'b000000;
12'b1011100011111: data = 6'b010101;
12'b1011100100000: data = 6'b010101;
12'b1011100100001: data = 6'b010101;
12'b1011100100010: data = 6'b010101;
12'b1011100100011: data = 6'b010101;
12'b1011100100100: data = 6'b010101;
12'b1011100100101: data = 6'b101001;
12'b1011100100110: data = 6'b101001;
12'b1011100100111: data = 6'b101010;
12'b1011100101000: data = 6'b101010;
12'b1011100101001: data = 6'b101010;
12'b1011100101010: data = 6'b101010;
12'b1011100101011: data = 6'b101010;
12'b1011100101100: data = 6'b101010;
12'b1011100101101: data = 6'b101010;
12'b1011100101110: data = 6'b101010;
12'b1011100101111: data = 6'b101010;
12'b1011100110000: data = 6'b101010;
12'b1011100110001: data = 6'b101010;
12'b1011100110010: data = 6'b101010;
12'b1011100110011: data = 6'b101010;
12'b1011100110100: data = 6'b101010;
12'b1011100110101: data = 6'b111010;
12'b1011100110110: data = 6'b111010;
12'b1011100110111: data = 6'b111110;
12'b1011100111000: data = 6'b111110;
12'b1011100111001: data = 6'b111111;
12'b1011100111010: data = 6'b111111;
12'b1011100111011: data = 6'b111111;
12'b1011100111100: data = 6'b111111;
12'b1011100111101: data = 6'b111111;
12'b1011100111110: data = 6'b111111;
12'b1011100111111: data = 6'b111111;
12'b10111001000000: data = 6'b111111;
12'b10111001000001: data = 6'b111111;
12'b10111001000010: data = 6'b111111;
12'b10111001000011: data = 6'b111111;
12'b10111001000100: data = 6'b111111;
12'b10111001000101: data = 6'b111111;
12'b10111001000110: data = 6'b111111;
12'b10111001000111: data = 6'b111110;
12'b10111001001000: data = 6'b111110;
12'b10111001001001: data = 6'b111110;
12'b10111001001010: data = 6'b111110;
12'b10111001001011: data = 6'b111110;
12'b10111001001100: data = 6'b111010;
12'b10111001001101: data = 6'b111010;
12'b10111001001110: data = 6'b111010;
12'b10111001001111: data = 6'b101010;
12'b10111001010000: data = 6'b101010;
12'b10111001010001: data = 6'b101010;
12'b10111001010010: data = 6'b101010;
12'b10111001010011: data = 6'b101010;
12'b10111001010100: data = 6'b101010;
12'b10111001010101: data = 6'b101010;
12'b10111001010110: data = 6'b101010;
12'b10111001010111: data = 6'b101010;
12'b10111001011000: data = 6'b101010;
12'b10111001011001: data = 6'b101010;
12'b10111001011010: data = 6'b101010;
12'b10111001011011: data = 6'b101010;
12'b10111001011100: data = 6'b101010;
12'b10111001011101: data = 6'b101010;
12'b10111001011110: data = 6'b101010;
12'b10111001011111: data = 6'b101010;
12'b10111001100000: data = 6'b101010;
12'b10111001100001: data = 6'b101010;
12'b10111001100010: data = 6'b101010;
12'b10111001100011: data = 6'b101010;
12'b10111001100100: data = 6'b101010;
12'b10111001100101: data = 6'b101010;
12'b10111001100110: data = 6'b101010;
12'b10111001100111: data = 6'b101010;
12'b10111001101000: data = 6'b101010;
12'b10111001101001: data = 6'b101010;
12'b10111001101010: data = 6'b101010;
12'b10111001101011: data = 6'b101010;
12'b10111001101100: data = 6'b101010;
12'b10111001101101: data = 6'b101010;
12'b10111001101110: data = 6'b101010;
12'b10111001101111: data = 6'b101010;
12'b10111001110000: data = 6'b101010;
12'b10111001110001: data = 6'b101010;
12'b10111001110010: data = 6'b101010;
12'b10111001110011: data = 6'b101010;
12'b10111001110100: data = 6'b101010;
12'b10111001110101: data = 6'b101010;
12'b10111001110110: data = 6'b101010;
12'b10111001110111: data = 6'b101010;
12'b10111001111000: data = 6'b101010;
12'b10111001111001: data = 6'b101001;
12'b10111001111010: data = 6'b101001;
12'b10111001111011: data = 6'b101001;
12'b10111001111100: data = 6'b010101;
12'b10111001111101: data = 6'b010101;
12'b10111001111110: data = 6'b010101;
12'b10111001111111: data = 6'b010101;
12'b101110010000000: data = 6'b010101;
12'b101110010000001: data = 6'b010101;
12'b101110010000010: data = 6'b010101;
12'b101110010000011: data = 6'b010101;
12'b101110010000100: data = 6'b010101;
12'b101110010000101: data = 6'b010101;
12'b101110010000110: data = 6'b010101;
12'b101110010000111: data = 6'b010101;
12'b101110010001000: data = 6'b010101;
12'b101110010001001: data = 6'b010101;
12'b101110010001010: data = 6'b010101;
12'b101110010001011: data = 6'b010101;
12'b101110010001100: data = 6'b000000;
12'b101110010001101: data = 6'b000000;
12'b101110010001110: data = 6'b101010;
12'b101110010001111: data = 6'b101010;
12'b101110010010000: data = 6'b101010;
12'b101110010010001: data = 6'b101010;
12'b101110010010010: data = 6'b010101;
12'b101110010010011: data = 6'b010101;
12'b101110010010100: data = 6'b010101;
12'b101110010010101: data = 6'b010101;
12'b101110010010110: data = 6'b010101;
12'b101110010010111: data = 6'b010101;
12'b101110010011000: data = 6'b010101;
12'b101110010011001: data = 6'b010101;
12'b101110010011010: data = 6'b010101;
12'b101110010011011: data = 6'b010101;
12'b101110010011100: data = 6'b010101;
12'b101110010011101: data = 6'b010101;
12'b101110010011110: data = 6'b010101;
12'b101110010011111: data = 6'b010101;
12'b101110010100000: data = 6'b010101;
12'b101110010100001: data = 6'b010101;
12'b101110010100010: data = 6'b010101;
12'b101110010100011: data = 6'b010101;
12'b101110010100100: data = 6'b010101;
12'b101110010100101: data = 6'b010101;
12'b101110010100110: data = 6'b010101;
12'b101110010100111: data = 6'b010101;
12'b101110010101000: data = 6'b010101;
12'b101110010101001: data = 6'b010101;
12'b101110010101010: data = 6'b010101;
12'b1011101000000: data = 6'b010101;
12'b1011101000001: data = 6'b010101;
12'b1011101000010: data = 6'b010101;
12'b1011101000011: data = 6'b010101;
12'b1011101000100: data = 6'b010101;
12'b1011101000101: data = 6'b010101;
12'b1011101000110: data = 6'b010101;
12'b1011101000111: data = 6'b010101;
12'b1011101001000: data = 6'b010101;
12'b1011101001001: data = 6'b010101;
12'b1011101001010: data = 6'b010101;
12'b1011101001011: data = 6'b010101;
12'b1011101001100: data = 6'b010101;
12'b1011101001101: data = 6'b010101;
12'b1011101001110: data = 6'b010101;
12'b1011101001111: data = 6'b010101;
12'b1011101010000: data = 6'b010101;
12'b1011101010001: data = 6'b010101;
12'b1011101010010: data = 6'b010101;
12'b1011101010011: data = 6'b010101;
12'b1011101010100: data = 6'b010101;
12'b1011101010101: data = 6'b010101;
12'b1011101010110: data = 6'b010101;
12'b1011101010111: data = 6'b010101;
12'b1011101011000: data = 6'b010101;
12'b1011101011001: data = 6'b101010;
12'b1011101011010: data = 6'b101010;
12'b1011101011011: data = 6'b101010;
12'b1011101011100: data = 6'b010101;
12'b1011101011101: data = 6'b000000;
12'b1011101011110: data = 6'b000000;
12'b1011101011111: data = 6'b010101;
12'b1011101100000: data = 6'b010101;
12'b1011101100001: data = 6'b010101;
12'b1011101100010: data = 6'b010101;
12'b1011101100011: data = 6'b010101;
12'b1011101100100: data = 6'b010101;
12'b1011101100101: data = 6'b101001;
12'b1011101100110: data = 6'b101001;
12'b1011101100111: data = 6'b101010;
12'b1011101101000: data = 6'b101010;
12'b1011101101001: data = 6'b101010;
12'b1011101101010: data = 6'b101010;
12'b1011101101011: data = 6'b101010;
12'b1011101101100: data = 6'b101010;
12'b1011101101101: data = 6'b101010;
12'b1011101101110: data = 6'b101010;
12'b1011101101111: data = 6'b101010;
12'b1011101110000: data = 6'b101010;
12'b1011101110001: data = 6'b101010;
12'b1011101110010: data = 6'b101010;
12'b1011101110011: data = 6'b101010;
12'b1011101110100: data = 6'b101010;
12'b1011101110101: data = 6'b111010;
12'b1011101110110: data = 6'b111010;
12'b1011101110111: data = 6'b111110;
12'b1011101111000: data = 6'b111110;
12'b1011101111001: data = 6'b111111;
12'b1011101111010: data = 6'b111111;
12'b1011101111011: data = 6'b111111;
12'b1011101111100: data = 6'b111111;
12'b1011101111101: data = 6'b111111;
12'b1011101111110: data = 6'b111111;
12'b1011101111111: data = 6'b111111;
12'b10111011000000: data = 6'b111111;
12'b10111011000001: data = 6'b111111;
12'b10111011000010: data = 6'b111111;
12'b10111011000011: data = 6'b111111;
12'b10111011000100: data = 6'b111111;
12'b10111011000101: data = 6'b111111;
12'b10111011000110: data = 6'b111111;
12'b10111011000111: data = 6'b111110;
12'b10111011001000: data = 6'b111110;
12'b10111011001001: data = 6'b111110;
12'b10111011001010: data = 6'b111110;
12'b10111011001011: data = 6'b111110;
12'b10111011001100: data = 6'b111010;
12'b10111011001101: data = 6'b111010;
12'b10111011001110: data = 6'b111010;
12'b10111011001111: data = 6'b101010;
12'b10111011010000: data = 6'b101010;
12'b10111011010001: data = 6'b101010;
12'b10111011010010: data = 6'b101010;
12'b10111011010011: data = 6'b101010;
12'b10111011010100: data = 6'b101010;
12'b10111011010101: data = 6'b101010;
12'b10111011010110: data = 6'b101010;
12'b10111011010111: data = 6'b101010;
12'b10111011011000: data = 6'b101010;
12'b10111011011001: data = 6'b101010;
12'b10111011011010: data = 6'b101010;
12'b10111011011011: data = 6'b101010;
12'b10111011011100: data = 6'b101010;
12'b10111011011101: data = 6'b101010;
12'b10111011011110: data = 6'b101010;
12'b10111011011111: data = 6'b101010;
12'b10111011100000: data = 6'b101010;
12'b10111011100001: data = 6'b101010;
12'b10111011100010: data = 6'b101010;
12'b10111011100011: data = 6'b101010;
12'b10111011100100: data = 6'b101010;
12'b10111011100101: data = 6'b101010;
12'b10111011100110: data = 6'b101010;
12'b10111011100111: data = 6'b101010;
12'b10111011101000: data = 6'b101010;
12'b10111011101001: data = 6'b101010;
12'b10111011101010: data = 6'b101010;
12'b10111011101011: data = 6'b101010;
12'b10111011101100: data = 6'b101010;
12'b10111011101101: data = 6'b101010;
12'b10111011101110: data = 6'b101010;
12'b10111011101111: data = 6'b101010;
12'b10111011110000: data = 6'b101010;
12'b10111011110001: data = 6'b101010;
12'b10111011110010: data = 6'b101010;
12'b10111011110011: data = 6'b101010;
12'b10111011110100: data = 6'b101010;
12'b10111011110101: data = 6'b101010;
12'b10111011110110: data = 6'b101010;
12'b10111011110111: data = 6'b101010;
12'b10111011111000: data = 6'b101010;
12'b10111011111001: data = 6'b101001;
12'b10111011111010: data = 6'b101001;
12'b10111011111011: data = 6'b101001;
12'b10111011111100: data = 6'b010101;
12'b10111011111101: data = 6'b010101;
12'b10111011111110: data = 6'b010101;
12'b10111011111111: data = 6'b010101;
12'b101110110000000: data = 6'b010101;
12'b101110110000001: data = 6'b010101;
12'b101110110000010: data = 6'b010101;
12'b101110110000011: data = 6'b010101;
12'b101110110000100: data = 6'b010101;
12'b101110110000101: data = 6'b010101;
12'b101110110000110: data = 6'b010101;
12'b101110110000111: data = 6'b010101;
12'b101110110001000: data = 6'b010101;
12'b101110110001001: data = 6'b010101;
12'b101110110001010: data = 6'b010101;
12'b101110110001011: data = 6'b010101;
12'b101110110001100: data = 6'b000000;
12'b101110110001101: data = 6'b000000;
12'b101110110001110: data = 6'b101010;
12'b101110110001111: data = 6'b101010;
12'b101110110010000: data = 6'b101010;
12'b101110110010001: data = 6'b101010;
12'b101110110010010: data = 6'b010101;
12'b101110110010011: data = 6'b010101;
12'b101110110010100: data = 6'b010101;
12'b101110110010101: data = 6'b010101;
12'b101110110010110: data = 6'b010101;
12'b101110110010111: data = 6'b010101;
12'b101110110011000: data = 6'b010101;
12'b101110110011001: data = 6'b010101;
12'b101110110011010: data = 6'b010101;
12'b101110110011011: data = 6'b010101;
12'b101110110011100: data = 6'b010101;
12'b101110110011101: data = 6'b010101;
12'b101110110011110: data = 6'b010101;
12'b101110110011111: data = 6'b010101;
12'b101110110100000: data = 6'b010101;
12'b101110110100001: data = 6'b010101;
12'b101110110100010: data = 6'b010101;
12'b101110110100011: data = 6'b010101;
12'b101110110100100: data = 6'b010101;
12'b101110110100101: data = 6'b010101;
12'b101110110100110: data = 6'b010101;
12'b101110110100111: data = 6'b010101;
12'b101110110101000: data = 6'b010101;
12'b101110110101001: data = 6'b010101;
12'b101110110101010: data = 6'b010101;
12'b1011110000000: data = 6'b010101;
12'b1011110000001: data = 6'b010101;
12'b1011110000010: data = 6'b010101;
12'b1011110000011: data = 6'b010101;
12'b1011110000100: data = 6'b010101;
12'b1011110000101: data = 6'b010101;
12'b1011110000110: data = 6'b010101;
12'b1011110000111: data = 6'b010101;
12'b1011110001000: data = 6'b010101;
12'b1011110001001: data = 6'b010101;
12'b1011110001010: data = 6'b010101;
12'b1011110001011: data = 6'b010101;
12'b1011110001100: data = 6'b010101;
12'b1011110001101: data = 6'b010101;
12'b1011110001110: data = 6'b010101;
12'b1011110001111: data = 6'b010101;
12'b1011110010000: data = 6'b010101;
12'b1011110010001: data = 6'b010101;
12'b1011110010010: data = 6'b010101;
12'b1011110010011: data = 6'b010101;
12'b1011110010100: data = 6'b010101;
12'b1011110010101: data = 6'b010101;
12'b1011110010110: data = 6'b010101;
12'b1011110010111: data = 6'b010101;
12'b1011110011000: data = 6'b010101;
12'b1011110011001: data = 6'b101010;
12'b1011110011010: data = 6'b101010;
12'b1011110011011: data = 6'b101010;
12'b1011110011100: data = 6'b010101;
12'b1011110011101: data = 6'b000000;
12'b1011110011110: data = 6'b000000;
12'b1011110011111: data = 6'b010101;
12'b1011110100000: data = 6'b010101;
12'b1011110100001: data = 6'b010101;
12'b1011110100010: data = 6'b010101;
12'b1011110100011: data = 6'b010101;
12'b1011110100100: data = 6'b010101;
12'b1011110100101: data = 6'b101001;
12'b1011110100110: data = 6'b101001;
12'b1011110100111: data = 6'b101010;
12'b1011110101000: data = 6'b101010;
12'b1011110101001: data = 6'b101010;
12'b1011110101010: data = 6'b101010;
12'b1011110101011: data = 6'b101010;
12'b1011110101100: data = 6'b101010;
12'b1011110101101: data = 6'b101010;
12'b1011110101110: data = 6'b101010;
12'b1011110101111: data = 6'b101010;
12'b1011110110000: data = 6'b101010;
12'b1011110110001: data = 6'b101010;
12'b1011110110010: data = 6'b101010;
12'b1011110110011: data = 6'b101010;
12'b1011110110100: data = 6'b101010;
12'b1011110110101: data = 6'b111010;
12'b1011110110110: data = 6'b111010;
12'b1011110110111: data = 6'b111110;
12'b1011110111000: data = 6'b111110;
12'b1011110111001: data = 6'b111111;
12'b1011110111010: data = 6'b111111;
12'b1011110111011: data = 6'b111111;
12'b1011110111100: data = 6'b111111;
12'b1011110111101: data = 6'b111111;
12'b1011110111110: data = 6'b111111;
12'b1011110111111: data = 6'b111111;
12'b10111101000000: data = 6'b111111;
12'b10111101000001: data = 6'b111111;
12'b10111101000010: data = 6'b111111;
12'b10111101000011: data = 6'b111111;
12'b10111101000100: data = 6'b111111;
12'b10111101000101: data = 6'b111111;
12'b10111101000110: data = 6'b111111;
12'b10111101000111: data = 6'b111110;
12'b10111101001000: data = 6'b111110;
12'b10111101001001: data = 6'b111110;
12'b10111101001010: data = 6'b111110;
12'b10111101001011: data = 6'b111110;
12'b10111101001100: data = 6'b111010;
12'b10111101001101: data = 6'b111010;
12'b10111101001110: data = 6'b111010;
12'b10111101001111: data = 6'b101010;
12'b10111101010000: data = 6'b101010;
12'b10111101010001: data = 6'b101010;
12'b10111101010010: data = 6'b101010;
12'b10111101010011: data = 6'b101010;
12'b10111101010100: data = 6'b101010;
12'b10111101010101: data = 6'b101010;
12'b10111101010110: data = 6'b101010;
12'b10111101010111: data = 6'b101010;
12'b10111101011000: data = 6'b101010;
12'b10111101011001: data = 6'b101010;
12'b10111101011010: data = 6'b101010;
12'b10111101011011: data = 6'b101010;
12'b10111101011100: data = 6'b101010;
12'b10111101011101: data = 6'b101010;
12'b10111101011110: data = 6'b101010;
12'b10111101011111: data = 6'b101010;
12'b10111101100000: data = 6'b101010;
12'b10111101100001: data = 6'b101010;
12'b10111101100010: data = 6'b101010;
12'b10111101100011: data = 6'b101010;
12'b10111101100100: data = 6'b101010;
12'b10111101100101: data = 6'b101010;
12'b10111101100110: data = 6'b101010;
12'b10111101100111: data = 6'b101010;
12'b10111101101000: data = 6'b101010;
12'b10111101101001: data = 6'b101010;
12'b10111101101010: data = 6'b101010;
12'b10111101101011: data = 6'b101010;
12'b10111101101100: data = 6'b101010;
12'b10111101101101: data = 6'b101010;
12'b10111101101110: data = 6'b101010;
12'b10111101101111: data = 6'b101010;
12'b10111101110000: data = 6'b101010;
12'b10111101110001: data = 6'b101010;
12'b10111101110010: data = 6'b101010;
12'b10111101110011: data = 6'b101010;
12'b10111101110100: data = 6'b101010;
12'b10111101110101: data = 6'b101010;
12'b10111101110110: data = 6'b101010;
12'b10111101110111: data = 6'b101010;
12'b10111101111000: data = 6'b101010;
12'b10111101111001: data = 6'b101001;
12'b10111101111010: data = 6'b101001;
12'b10111101111011: data = 6'b101001;
12'b10111101111100: data = 6'b010101;
12'b10111101111101: data = 6'b010101;
12'b10111101111110: data = 6'b010101;
12'b10111101111111: data = 6'b010101;
12'b101111010000000: data = 6'b010101;
12'b101111010000001: data = 6'b010101;
12'b101111010000010: data = 6'b010101;
12'b101111010000011: data = 6'b010101;
12'b101111010000100: data = 6'b010101;
12'b101111010000101: data = 6'b010101;
12'b101111010000110: data = 6'b010101;
12'b101111010000111: data = 6'b010101;
12'b101111010001000: data = 6'b010101;
12'b101111010001001: data = 6'b010101;
12'b101111010001010: data = 6'b010101;
12'b101111010001011: data = 6'b010101;
12'b101111010001100: data = 6'b000000;
12'b101111010001101: data = 6'b000000;
12'b101111010001110: data = 6'b101010;
12'b101111010001111: data = 6'b101010;
12'b101111010010000: data = 6'b101010;
12'b101111010010001: data = 6'b101010;
12'b101111010010010: data = 6'b010101;
12'b101111010010011: data = 6'b010101;
12'b101111010010100: data = 6'b010101;
12'b101111010010101: data = 6'b010101;
12'b101111010010110: data = 6'b010101;
12'b101111010010111: data = 6'b010101;
12'b101111010011000: data = 6'b010101;
12'b101111010011001: data = 6'b010101;
12'b101111010011010: data = 6'b010101;
12'b101111010011011: data = 6'b010101;
12'b101111010011100: data = 6'b010101;
12'b101111010011101: data = 6'b010101;
12'b101111010011110: data = 6'b010101;
12'b101111010011111: data = 6'b010101;
12'b101111010100000: data = 6'b010101;
12'b101111010100001: data = 6'b010101;
12'b101111010100010: data = 6'b010101;
12'b101111010100011: data = 6'b010101;
12'b101111010100100: data = 6'b010101;
12'b101111010100101: data = 6'b010101;
12'b101111010100110: data = 6'b010101;
12'b101111010100111: data = 6'b010101;
12'b101111010101000: data = 6'b010101;
12'b101111010101001: data = 6'b010101;
12'b101111010101010: data = 6'b010101;
12'b1011111000000: data = 6'b010101;
12'b1011111000001: data = 6'b010101;
12'b1011111000010: data = 6'b010101;
12'b1011111000011: data = 6'b010101;
12'b1011111000100: data = 6'b010101;
12'b1011111000101: data = 6'b010101;
12'b1011111000110: data = 6'b010101;
12'b1011111000111: data = 6'b010101;
12'b1011111001000: data = 6'b010101;
12'b1011111001001: data = 6'b010101;
12'b1011111001010: data = 6'b010101;
12'b1011111001011: data = 6'b010101;
12'b1011111001100: data = 6'b010101;
12'b1011111001101: data = 6'b010101;
12'b1011111001110: data = 6'b010101;
12'b1011111001111: data = 6'b010101;
12'b1011111010000: data = 6'b010101;
12'b1011111010001: data = 6'b010101;
12'b1011111010010: data = 6'b010101;
12'b1011111010011: data = 6'b010101;
12'b1011111010100: data = 6'b010101;
12'b1011111010101: data = 6'b010101;
12'b1011111010110: data = 6'b010101;
12'b1011111010111: data = 6'b010101;
12'b1011111011000: data = 6'b010101;
12'b1011111011001: data = 6'b101010;
12'b1011111011010: data = 6'b101010;
12'b1011111011011: data = 6'b101010;
12'b1011111011100: data = 6'b010101;
12'b1011111011101: data = 6'b000000;
12'b1011111011110: data = 6'b000000;
12'b1011111011111: data = 6'b010101;
12'b1011111100000: data = 6'b010101;
12'b1011111100001: data = 6'b010101;
12'b1011111100010: data = 6'b010101;
12'b1011111100011: data = 6'b010101;
12'b1011111100100: data = 6'b010101;
12'b1011111100101: data = 6'b101001;
12'b1011111100110: data = 6'b101001;
12'b1011111100111: data = 6'b101010;
12'b1011111101000: data = 6'b101010;
12'b1011111101001: data = 6'b101010;
12'b1011111101010: data = 6'b101010;
12'b1011111101011: data = 6'b101010;
12'b1011111101100: data = 6'b101010;
12'b1011111101101: data = 6'b101010;
12'b1011111101110: data = 6'b101010;
12'b1011111101111: data = 6'b101010;
12'b1011111110000: data = 6'b101010;
12'b1011111110001: data = 6'b101010;
12'b1011111110010: data = 6'b101010;
12'b1011111110011: data = 6'b101010;
12'b1011111110100: data = 6'b101010;
12'b1011111110101: data = 6'b111010;
12'b1011111110110: data = 6'b111010;
12'b1011111110111: data = 6'b111110;
12'b1011111111000: data = 6'b111110;
12'b1011111111001: data = 6'b111111;
12'b1011111111010: data = 6'b111111;
12'b1011111111011: data = 6'b111111;
12'b1011111111100: data = 6'b111111;
12'b1011111111101: data = 6'b111111;
12'b1011111111110: data = 6'b111111;
12'b1011111111111: data = 6'b111111;
12'b10111111000000: data = 6'b111111;
12'b10111111000001: data = 6'b111111;
12'b10111111000010: data = 6'b111111;
12'b10111111000011: data = 6'b111111;
12'b10111111000100: data = 6'b111111;
12'b10111111000101: data = 6'b111111;
12'b10111111000110: data = 6'b111111;
12'b10111111000111: data = 6'b111110;
12'b10111111001000: data = 6'b111110;
12'b10111111001001: data = 6'b111110;
12'b10111111001010: data = 6'b111110;
12'b10111111001011: data = 6'b111110;
12'b10111111001100: data = 6'b111010;
12'b10111111001101: data = 6'b111010;
12'b10111111001110: data = 6'b111010;
12'b10111111001111: data = 6'b101010;
12'b10111111010000: data = 6'b101010;
12'b10111111010001: data = 6'b101010;
12'b10111111010010: data = 6'b101010;
12'b10111111010011: data = 6'b101010;
12'b10111111010100: data = 6'b101010;
12'b10111111010101: data = 6'b101010;
12'b10111111010110: data = 6'b101010;
12'b10111111010111: data = 6'b101010;
12'b10111111011000: data = 6'b101010;
12'b10111111011001: data = 6'b101010;
12'b10111111011010: data = 6'b101010;
12'b10111111011011: data = 6'b101010;
12'b10111111011100: data = 6'b101010;
12'b10111111011101: data = 6'b101010;
12'b10111111011110: data = 6'b101010;
12'b10111111011111: data = 6'b101010;
12'b10111111100000: data = 6'b101010;
12'b10111111100001: data = 6'b101010;
12'b10111111100010: data = 6'b101010;
12'b10111111100011: data = 6'b101010;
12'b10111111100100: data = 6'b101010;
12'b10111111100101: data = 6'b101010;
12'b10111111100110: data = 6'b101010;
12'b10111111100111: data = 6'b101010;
12'b10111111101000: data = 6'b101010;
12'b10111111101001: data = 6'b101010;
12'b10111111101010: data = 6'b101010;
12'b10111111101011: data = 6'b101010;
12'b10111111101100: data = 6'b101010;
12'b10111111101101: data = 6'b101010;
12'b10111111101110: data = 6'b101010;
12'b10111111101111: data = 6'b101010;
12'b10111111110000: data = 6'b101010;
12'b10111111110001: data = 6'b101010;
12'b10111111110010: data = 6'b101010;
12'b10111111110011: data = 6'b101010;
12'b10111111110100: data = 6'b101010;
12'b10111111110101: data = 6'b101010;
12'b10111111110110: data = 6'b101010;
12'b10111111110111: data = 6'b101010;
12'b10111111111000: data = 6'b101010;
12'b10111111111001: data = 6'b101001;
12'b10111111111010: data = 6'b101001;
12'b10111111111011: data = 6'b101001;
12'b10111111111100: data = 6'b010101;
12'b10111111111101: data = 6'b010101;
12'b10111111111110: data = 6'b010101;
12'b10111111111111: data = 6'b010101;
12'b101111110000000: data = 6'b010101;
12'b101111110000001: data = 6'b010101;
12'b101111110000010: data = 6'b010101;
12'b101111110000011: data = 6'b010101;
12'b101111110000100: data = 6'b010101;
12'b101111110000101: data = 6'b010101;
12'b101111110000110: data = 6'b010101;
12'b101111110000111: data = 6'b010101;
12'b101111110001000: data = 6'b010101;
12'b101111110001001: data = 6'b010101;
12'b101111110001010: data = 6'b010101;
12'b101111110001011: data = 6'b010101;
12'b101111110001100: data = 6'b000000;
12'b101111110001101: data = 6'b000000;
12'b101111110001110: data = 6'b101010;
12'b101111110001111: data = 6'b101010;
12'b101111110010000: data = 6'b101010;
12'b101111110010001: data = 6'b101010;
12'b101111110010010: data = 6'b010101;
12'b101111110010011: data = 6'b010101;
12'b101111110010100: data = 6'b010101;
12'b101111110010101: data = 6'b010101;
12'b101111110010110: data = 6'b010101;
12'b101111110010111: data = 6'b010101;
12'b101111110011000: data = 6'b010101;
12'b101111110011001: data = 6'b010101;
12'b101111110011010: data = 6'b010101;
12'b101111110011011: data = 6'b010101;
12'b101111110011100: data = 6'b010101;
12'b101111110011101: data = 6'b010101;
12'b101111110011110: data = 6'b010101;
12'b101111110011111: data = 6'b010101;
12'b101111110100000: data = 6'b010101;
12'b101111110100001: data = 6'b010101;
12'b101111110100010: data = 6'b010101;
12'b101111110100011: data = 6'b010101;
12'b101111110100100: data = 6'b010101;
12'b101111110100101: data = 6'b010101;
12'b101111110100110: data = 6'b010101;
12'b101111110100111: data = 6'b010101;
12'b101111110101000: data = 6'b010101;
12'b101111110101001: data = 6'b010101;
12'b101111110101010: data = 6'b010101;
12'b1100000000000: data = 6'b010101;
12'b1100000000001: data = 6'b010101;
12'b1100000000010: data = 6'b010101;
12'b1100000000011: data = 6'b010101;
12'b1100000000100: data = 6'b010101;
12'b1100000000101: data = 6'b010101;
12'b1100000000110: data = 6'b010101;
12'b1100000000111: data = 6'b010101;
12'b1100000001000: data = 6'b010101;
12'b1100000001001: data = 6'b010101;
12'b1100000001010: data = 6'b010101;
12'b1100000001011: data = 6'b010101;
12'b1100000001100: data = 6'b010101;
12'b1100000001101: data = 6'b010101;
12'b1100000001110: data = 6'b010101;
12'b1100000001111: data = 6'b010101;
12'b1100000010000: data = 6'b010101;
12'b1100000010001: data = 6'b010101;
12'b1100000010010: data = 6'b010101;
12'b1100000010011: data = 6'b010101;
12'b1100000010100: data = 6'b010101;
12'b1100000010101: data = 6'b010101;
12'b1100000010110: data = 6'b010101;
12'b1100000010111: data = 6'b010101;
12'b1100000011000: data = 6'b010101;
12'b1100000011001: data = 6'b101010;
12'b1100000011010: data = 6'b101010;
12'b1100000011011: data = 6'b101010;
12'b1100000011100: data = 6'b010101;
12'b1100000011101: data = 6'b000000;
12'b1100000011110: data = 6'b000000;
12'b1100000011111: data = 6'b010101;
12'b1100000100000: data = 6'b010101;
12'b1100000100001: data = 6'b010101;
12'b1100000100010: data = 6'b010101;
12'b1100000100011: data = 6'b010101;
12'b1100000100100: data = 6'b010101;
12'b1100000100101: data = 6'b101001;
12'b1100000100110: data = 6'b101001;
12'b1100000100111: data = 6'b101010;
12'b1100000101000: data = 6'b101010;
12'b1100000101001: data = 6'b101010;
12'b1100000101010: data = 6'b101010;
12'b1100000101011: data = 6'b101010;
12'b1100000101100: data = 6'b101010;
12'b1100000101101: data = 6'b101010;
12'b1100000101110: data = 6'b101010;
12'b1100000101111: data = 6'b101010;
12'b1100000110000: data = 6'b101010;
12'b1100000110001: data = 6'b101010;
12'b1100000110010: data = 6'b101010;
12'b1100000110011: data = 6'b101010;
12'b1100000110100: data = 6'b101010;
12'b1100000110101: data = 6'b111010;
12'b1100000110110: data = 6'b111010;
12'b1100000110111: data = 6'b111110;
12'b1100000111000: data = 6'b111110;
12'b1100000111001: data = 6'b111111;
12'b1100000111010: data = 6'b111111;
12'b1100000111011: data = 6'b111111;
12'b1100000111100: data = 6'b111111;
12'b1100000111101: data = 6'b111111;
12'b1100000111110: data = 6'b111111;
12'b1100000111111: data = 6'b111111;
12'b11000001000000: data = 6'b111111;
12'b11000001000001: data = 6'b111111;
12'b11000001000010: data = 6'b111111;
12'b11000001000011: data = 6'b111111;
12'b11000001000100: data = 6'b111111;
12'b11000001000101: data = 6'b111111;
12'b11000001000110: data = 6'b111111;
12'b11000001000111: data = 6'b111110;
12'b11000001001000: data = 6'b111110;
12'b11000001001001: data = 6'b111110;
12'b11000001001010: data = 6'b111110;
12'b11000001001011: data = 6'b111110;
12'b11000001001100: data = 6'b111010;
12'b11000001001101: data = 6'b111010;
12'b11000001001110: data = 6'b101010;
12'b11000001001111: data = 6'b101010;
12'b11000001010000: data = 6'b101010;
12'b11000001010001: data = 6'b101010;
12'b11000001010010: data = 6'b101010;
12'b11000001010011: data = 6'b101010;
12'b11000001010100: data = 6'b101010;
12'b11000001010101: data = 6'b101010;
12'b11000001010110: data = 6'b101010;
12'b11000001010111: data = 6'b101010;
12'b11000001011000: data = 6'b101010;
12'b11000001011001: data = 6'b101010;
12'b11000001011010: data = 6'b101010;
12'b11000001011011: data = 6'b101010;
12'b11000001011100: data = 6'b101010;
12'b11000001011101: data = 6'b101010;
12'b11000001011110: data = 6'b101010;
12'b11000001011111: data = 6'b101010;
12'b11000001100000: data = 6'b101010;
12'b11000001100001: data = 6'b101010;
12'b11000001100010: data = 6'b101010;
12'b11000001100011: data = 6'b101010;
12'b11000001100100: data = 6'b101010;
12'b11000001100101: data = 6'b101010;
12'b11000001100110: data = 6'b101010;
12'b11000001100111: data = 6'b101010;
12'b11000001101000: data = 6'b101010;
12'b11000001101001: data = 6'b101010;
12'b11000001101010: data = 6'b101010;
12'b11000001101011: data = 6'b101010;
12'b11000001101100: data = 6'b101010;
12'b11000001101101: data = 6'b101010;
12'b11000001101110: data = 6'b101010;
12'b11000001101111: data = 6'b101010;
12'b11000001110000: data = 6'b101010;
12'b11000001110001: data = 6'b101010;
12'b11000001110010: data = 6'b101010;
12'b11000001110011: data = 6'b101010;
12'b11000001110100: data = 6'b101010;
12'b11000001110101: data = 6'b101010;
12'b11000001110110: data = 6'b101010;
12'b11000001110111: data = 6'b101010;
12'b11000001111000: data = 6'b101010;
12'b11000001111001: data = 6'b101001;
12'b11000001111010: data = 6'b101001;
12'b11000001111011: data = 6'b101001;
12'b11000001111100: data = 6'b010101;
12'b11000001111101: data = 6'b010101;
12'b11000001111110: data = 6'b010101;
12'b11000001111111: data = 6'b010101;
12'b110000010000000: data = 6'b010101;
12'b110000010000001: data = 6'b010101;
12'b110000010000010: data = 6'b010101;
12'b110000010000011: data = 6'b010101;
12'b110000010000100: data = 6'b010101;
12'b110000010000101: data = 6'b010101;
12'b110000010000110: data = 6'b010101;
12'b110000010000111: data = 6'b010101;
12'b110000010001000: data = 6'b010101;
12'b110000010001001: data = 6'b010101;
12'b110000010001010: data = 6'b010101;
12'b110000010001011: data = 6'b010101;
12'b110000010001100: data = 6'b000000;
12'b110000010001101: data = 6'b000000;
12'b110000010001110: data = 6'b101010;
12'b110000010001111: data = 6'b101010;
12'b110000010010000: data = 6'b101010;
12'b110000010010001: data = 6'b101010;
12'b110000010010010: data = 6'b010101;
12'b110000010010011: data = 6'b010101;
12'b110000010010100: data = 6'b010101;
12'b110000010010101: data = 6'b010101;
12'b110000010010110: data = 6'b010101;
12'b110000010010111: data = 6'b010101;
12'b110000010011000: data = 6'b010101;
12'b110000010011001: data = 6'b010101;
12'b110000010011010: data = 6'b010101;
12'b110000010011011: data = 6'b010101;
12'b110000010011100: data = 6'b010101;
12'b110000010011101: data = 6'b010101;
12'b110000010011110: data = 6'b010101;
12'b110000010011111: data = 6'b010101;
12'b110000010100000: data = 6'b010101;
12'b110000010100001: data = 6'b010101;
12'b110000010100010: data = 6'b010101;
12'b110000010100011: data = 6'b010101;
12'b110000010100100: data = 6'b010101;
12'b110000010100101: data = 6'b010101;
12'b110000010100110: data = 6'b010101;
12'b110000010100111: data = 6'b010101;
12'b110000010101000: data = 6'b010101;
12'b110000010101001: data = 6'b010101;
12'b110000010101010: data = 6'b010101;
12'b1100001000000: data = 6'b010101;
12'b1100001000001: data = 6'b010101;
12'b1100001000010: data = 6'b010101;
12'b1100001000011: data = 6'b010101;
12'b1100001000100: data = 6'b010101;
12'b1100001000101: data = 6'b010101;
12'b1100001000110: data = 6'b010101;
12'b1100001000111: data = 6'b010101;
12'b1100001001000: data = 6'b010101;
12'b1100001001001: data = 6'b010101;
12'b1100001001010: data = 6'b010101;
12'b1100001001011: data = 6'b010101;
12'b1100001001100: data = 6'b010101;
12'b1100001001101: data = 6'b010101;
12'b1100001001110: data = 6'b010101;
12'b1100001001111: data = 6'b010101;
12'b1100001010000: data = 6'b010101;
12'b1100001010001: data = 6'b010101;
12'b1100001010010: data = 6'b010101;
12'b1100001010011: data = 6'b010101;
12'b1100001010100: data = 6'b010101;
12'b1100001010101: data = 6'b010101;
12'b1100001010110: data = 6'b010101;
12'b1100001010111: data = 6'b010101;
12'b1100001011000: data = 6'b010101;
12'b1100001011001: data = 6'b101010;
12'b1100001011010: data = 6'b101010;
12'b1100001011011: data = 6'b101010;
12'b1100001011100: data = 6'b010101;
12'b1100001011101: data = 6'b000000;
12'b1100001011110: data = 6'b000000;
12'b1100001011111: data = 6'b010101;
12'b1100001100000: data = 6'b010101;
12'b1100001100001: data = 6'b010101;
12'b1100001100010: data = 6'b010101;
12'b1100001100011: data = 6'b010101;
12'b1100001100100: data = 6'b010101;
12'b1100001100101: data = 6'b101001;
12'b1100001100110: data = 6'b101001;
12'b1100001100111: data = 6'b101010;
12'b1100001101000: data = 6'b101010;
12'b1100001101001: data = 6'b101010;
12'b1100001101010: data = 6'b101010;
12'b1100001101011: data = 6'b101010;
12'b1100001101100: data = 6'b101010;
12'b1100001101101: data = 6'b101010;
12'b1100001101110: data = 6'b101010;
12'b1100001101111: data = 6'b101010;
12'b1100001110000: data = 6'b101010;
12'b1100001110001: data = 6'b101010;
12'b1100001110010: data = 6'b101010;
12'b1100001110011: data = 6'b101010;
12'b1100001110100: data = 6'b101010;
12'b1100001110101: data = 6'b111010;
12'b1100001110110: data = 6'b111010;
12'b1100001110111: data = 6'b111110;
12'b1100001111000: data = 6'b111110;
12'b1100001111001: data = 6'b111111;
12'b1100001111010: data = 6'b111111;
12'b1100001111011: data = 6'b111111;
12'b1100001111100: data = 6'b111111;
12'b1100001111101: data = 6'b111111;
12'b1100001111110: data = 6'b111111;
12'b1100001111111: data = 6'b111111;
12'b11000011000000: data = 6'b111111;
12'b11000011000001: data = 6'b111111;
12'b11000011000010: data = 6'b111111;
12'b11000011000011: data = 6'b111111;
12'b11000011000100: data = 6'b111111;
12'b11000011000101: data = 6'b111111;
12'b11000011000110: data = 6'b111111;
12'b11000011000111: data = 6'b111110;
12'b11000011001000: data = 6'b111110;
12'b11000011001001: data = 6'b111110;
12'b11000011001010: data = 6'b111110;
12'b11000011001011: data = 6'b111110;
12'b11000011001100: data = 6'b111010;
12'b11000011001101: data = 6'b111010;
12'b11000011001110: data = 6'b111010;
12'b11000011001111: data = 6'b101010;
12'b11000011010000: data = 6'b101010;
12'b11000011010001: data = 6'b101010;
12'b11000011010010: data = 6'b101010;
12'b11000011010011: data = 6'b101010;
12'b11000011010100: data = 6'b101010;
12'b11000011010101: data = 6'b101010;
12'b11000011010110: data = 6'b101010;
12'b11000011010111: data = 6'b101010;
12'b11000011011000: data = 6'b101010;
12'b11000011011001: data = 6'b101010;
12'b11000011011010: data = 6'b101010;
12'b11000011011011: data = 6'b101010;
12'b11000011011100: data = 6'b101010;
12'b11000011011101: data = 6'b101010;
12'b11000011011110: data = 6'b101010;
12'b11000011011111: data = 6'b101010;
12'b11000011100000: data = 6'b101010;
12'b11000011100001: data = 6'b101010;
12'b11000011100010: data = 6'b101010;
12'b11000011100011: data = 6'b101010;
12'b11000011100100: data = 6'b101010;
12'b11000011100101: data = 6'b101010;
12'b11000011100110: data = 6'b101010;
12'b11000011100111: data = 6'b101010;
12'b11000011101000: data = 6'b101010;
12'b11000011101001: data = 6'b101010;
12'b11000011101010: data = 6'b101010;
12'b11000011101011: data = 6'b101010;
12'b11000011101100: data = 6'b101010;
12'b11000011101101: data = 6'b101010;
12'b11000011101110: data = 6'b101010;
12'b11000011101111: data = 6'b101010;
12'b11000011110000: data = 6'b101010;
12'b11000011110001: data = 6'b101010;
12'b11000011110010: data = 6'b101010;
12'b11000011110011: data = 6'b101010;
12'b11000011110100: data = 6'b101010;
12'b11000011110101: data = 6'b101010;
12'b11000011110110: data = 6'b101010;
12'b11000011110111: data = 6'b101010;
12'b11000011111000: data = 6'b101010;
12'b11000011111001: data = 6'b101001;
12'b11000011111010: data = 6'b101001;
12'b11000011111011: data = 6'b101001;
12'b11000011111100: data = 6'b010101;
12'b11000011111101: data = 6'b010101;
12'b11000011111110: data = 6'b010101;
12'b11000011111111: data = 6'b010101;
12'b110000110000000: data = 6'b010101;
12'b110000110000001: data = 6'b010101;
12'b110000110000010: data = 6'b010101;
12'b110000110000011: data = 6'b010101;
12'b110000110000100: data = 6'b010101;
12'b110000110000101: data = 6'b010101;
12'b110000110000110: data = 6'b010101;
12'b110000110000111: data = 6'b010101;
12'b110000110001000: data = 6'b010101;
12'b110000110001001: data = 6'b010101;
12'b110000110001010: data = 6'b010101;
12'b110000110001011: data = 6'b010101;
12'b110000110001100: data = 6'b000000;
12'b110000110001101: data = 6'b000000;
12'b110000110001110: data = 6'b101010;
12'b110000110001111: data = 6'b101010;
12'b110000110010000: data = 6'b101010;
12'b110000110010001: data = 6'b101010;
12'b110000110010010: data = 6'b010101;
12'b110000110010011: data = 6'b010101;
12'b110000110010100: data = 6'b010101;
12'b110000110010101: data = 6'b010101;
12'b110000110010110: data = 6'b010101;
12'b110000110010111: data = 6'b010101;
12'b110000110011000: data = 6'b010101;
12'b110000110011001: data = 6'b010101;
12'b110000110011010: data = 6'b010101;
12'b110000110011011: data = 6'b010101;
12'b110000110011100: data = 6'b010101;
12'b110000110011101: data = 6'b010101;
12'b110000110011110: data = 6'b010101;
12'b110000110011111: data = 6'b010101;
12'b110000110100000: data = 6'b010101;
12'b110000110100001: data = 6'b010101;
12'b110000110100010: data = 6'b010101;
12'b110000110100011: data = 6'b010101;
12'b110000110100100: data = 6'b010101;
12'b110000110100101: data = 6'b010101;
12'b110000110100110: data = 6'b010101;
12'b110000110100111: data = 6'b010101;
12'b110000110101000: data = 6'b010101;
12'b110000110101001: data = 6'b010101;
12'b110000110101010: data = 6'b010101;
12'b1100010000000: data = 6'b010101;
12'b1100010000001: data = 6'b010101;
12'b1100010000010: data = 6'b010101;
12'b1100010000011: data = 6'b010101;
12'b1100010000100: data = 6'b010101;
12'b1100010000101: data = 6'b010101;
12'b1100010000110: data = 6'b010101;
12'b1100010000111: data = 6'b010101;
12'b1100010001000: data = 6'b010101;
12'b1100010001001: data = 6'b010101;
12'b1100010001010: data = 6'b010101;
12'b1100010001011: data = 6'b010101;
12'b1100010001100: data = 6'b010101;
12'b1100010001101: data = 6'b010101;
12'b1100010001110: data = 6'b010101;
12'b1100010001111: data = 6'b010101;
12'b1100010010000: data = 6'b010101;
12'b1100010010001: data = 6'b010101;
12'b1100010010010: data = 6'b010101;
12'b1100010010011: data = 6'b010101;
12'b1100010010100: data = 6'b010101;
12'b1100010010101: data = 6'b010101;
12'b1100010010110: data = 6'b010101;
12'b1100010010111: data = 6'b010101;
12'b1100010011000: data = 6'b010101;
12'b1100010011001: data = 6'b101010;
12'b1100010011010: data = 6'b101010;
12'b1100010011011: data = 6'b101010;
12'b1100010011100: data = 6'b010101;
12'b1100010011101: data = 6'b000000;
12'b1100010011110: data = 6'b000000;
12'b1100010011111: data = 6'b010101;
12'b1100010100000: data = 6'b010101;
12'b1100010100001: data = 6'b010101;
12'b1100010100010: data = 6'b010101;
12'b1100010100011: data = 6'b010101;
12'b1100010100100: data = 6'b010101;
12'b1100010100101: data = 6'b101001;
12'b1100010100110: data = 6'b101001;
12'b1100010100111: data = 6'b101010;
12'b1100010101000: data = 6'b101010;
12'b1100010101001: data = 6'b101010;
12'b1100010101010: data = 6'b101010;
12'b1100010101011: data = 6'b101010;
12'b1100010101100: data = 6'b101010;
12'b1100010101101: data = 6'b101010;
12'b1100010101110: data = 6'b101010;
12'b1100010101111: data = 6'b101010;
12'b1100010110000: data = 6'b101010;
12'b1100010110001: data = 6'b101010;
12'b1100010110010: data = 6'b101010;
12'b1100010110011: data = 6'b101010;
12'b1100010110100: data = 6'b101010;
12'b1100010110101: data = 6'b111010;
12'b1100010110110: data = 6'b111010;
12'b1100010110111: data = 6'b111110;
12'b1100010111000: data = 6'b111110;
12'b1100010111001: data = 6'b111111;
12'b1100010111010: data = 6'b111111;
12'b1100010111011: data = 6'b111111;
12'b1100010111100: data = 6'b111111;
12'b1100010111101: data = 6'b111111;
12'b1100010111110: data = 6'b111111;
12'b1100010111111: data = 6'b111111;
12'b11000101000000: data = 6'b111111;
12'b11000101000001: data = 6'b111111;
12'b11000101000010: data = 6'b111111;
12'b11000101000011: data = 6'b111111;
12'b11000101000100: data = 6'b111111;
12'b11000101000101: data = 6'b111111;
12'b11000101000110: data = 6'b111111;
12'b11000101000111: data = 6'b111110;
12'b11000101001000: data = 6'b111110;
12'b11000101001001: data = 6'b111110;
12'b11000101001010: data = 6'b111110;
12'b11000101001011: data = 6'b111110;
12'b11000101001100: data = 6'b111010;
12'b11000101001101: data = 6'b111010;
12'b11000101001110: data = 6'b101010;
12'b11000101001111: data = 6'b101010;
12'b11000101010000: data = 6'b101010;
12'b11000101010001: data = 6'b101010;
12'b11000101010010: data = 6'b101010;
12'b11000101010011: data = 6'b101010;
12'b11000101010100: data = 6'b101010;
12'b11000101010101: data = 6'b101010;
12'b11000101010110: data = 6'b101010;
12'b11000101010111: data = 6'b101010;
12'b11000101011000: data = 6'b101010;
12'b11000101011001: data = 6'b101010;
12'b11000101011010: data = 6'b101010;
12'b11000101011011: data = 6'b101010;
12'b11000101011100: data = 6'b101010;
12'b11000101011101: data = 6'b101010;
12'b11000101011110: data = 6'b101010;
12'b11000101011111: data = 6'b101010;
12'b11000101100000: data = 6'b101010;
12'b11000101100001: data = 6'b101010;
12'b11000101100010: data = 6'b101010;
12'b11000101100011: data = 6'b101010;
12'b11000101100100: data = 6'b101010;
12'b11000101100101: data = 6'b101010;
12'b11000101100110: data = 6'b101010;
12'b11000101100111: data = 6'b101010;
12'b11000101101000: data = 6'b101010;
12'b11000101101001: data = 6'b101010;
12'b11000101101010: data = 6'b101010;
12'b11000101101011: data = 6'b101010;
12'b11000101101100: data = 6'b101010;
12'b11000101101101: data = 6'b101010;
12'b11000101101110: data = 6'b101010;
12'b11000101101111: data = 6'b101010;
12'b11000101110000: data = 6'b101010;
12'b11000101110001: data = 6'b101010;
12'b11000101110010: data = 6'b101010;
12'b11000101110011: data = 6'b101010;
12'b11000101110100: data = 6'b101010;
12'b11000101110101: data = 6'b101010;
12'b11000101110110: data = 6'b101010;
12'b11000101110111: data = 6'b101010;
12'b11000101111000: data = 6'b101010;
12'b11000101111001: data = 6'b101001;
12'b11000101111010: data = 6'b101001;
12'b11000101111011: data = 6'b101001;
12'b11000101111100: data = 6'b010101;
12'b11000101111101: data = 6'b010101;
12'b11000101111110: data = 6'b010101;
12'b11000101111111: data = 6'b010101;
12'b110001010000000: data = 6'b010101;
12'b110001010000001: data = 6'b010101;
12'b110001010000010: data = 6'b010101;
12'b110001010000011: data = 6'b010101;
12'b110001010000100: data = 6'b010101;
12'b110001010000101: data = 6'b010101;
12'b110001010000110: data = 6'b010101;
12'b110001010000111: data = 6'b010101;
12'b110001010001000: data = 6'b010101;
12'b110001010001001: data = 6'b010101;
12'b110001010001010: data = 6'b010101;
12'b110001010001011: data = 6'b010101;
12'b110001010001100: data = 6'b000000;
12'b110001010001101: data = 6'b000000;
12'b110001010001110: data = 6'b101010;
12'b110001010001111: data = 6'b101010;
12'b110001010010000: data = 6'b101010;
12'b110001010010001: data = 6'b101010;
12'b110001010010010: data = 6'b010101;
12'b110001010010011: data = 6'b010101;
12'b110001010010100: data = 6'b010101;
12'b110001010010101: data = 6'b010101;
12'b110001010010110: data = 6'b010101;
12'b110001010010111: data = 6'b010101;
12'b110001010011000: data = 6'b010101;
12'b110001010011001: data = 6'b010101;
12'b110001010011010: data = 6'b010101;
12'b110001010011011: data = 6'b010101;
12'b110001010011100: data = 6'b010101;
12'b110001010011101: data = 6'b010101;
12'b110001010011110: data = 6'b010101;
12'b110001010011111: data = 6'b010101;
12'b110001010100000: data = 6'b010101;
12'b110001010100001: data = 6'b010101;
12'b110001010100010: data = 6'b010101;
12'b110001010100011: data = 6'b010101;
12'b110001010100100: data = 6'b010101;
12'b110001010100101: data = 6'b010101;
12'b110001010100110: data = 6'b010101;
12'b110001010100111: data = 6'b010101;
12'b110001010101000: data = 6'b010101;
12'b110001010101001: data = 6'b010101;
12'b110001010101010: data = 6'b010101;
12'b1100011000000: data = 6'b010101;
12'b1100011000001: data = 6'b010101;
12'b1100011000010: data = 6'b010101;
12'b1100011000011: data = 6'b010101;
12'b1100011000100: data = 6'b010101;
12'b1100011000101: data = 6'b010101;
12'b1100011000110: data = 6'b010101;
12'b1100011000111: data = 6'b010101;
12'b1100011001000: data = 6'b010101;
12'b1100011001001: data = 6'b010101;
12'b1100011001010: data = 6'b010101;
12'b1100011001011: data = 6'b010101;
12'b1100011001100: data = 6'b010101;
12'b1100011001101: data = 6'b010101;
12'b1100011001110: data = 6'b010101;
12'b1100011001111: data = 6'b010101;
12'b1100011010000: data = 6'b010101;
12'b1100011010001: data = 6'b010101;
12'b1100011010010: data = 6'b010101;
12'b1100011010011: data = 6'b010101;
12'b1100011010100: data = 6'b010101;
12'b1100011010101: data = 6'b010101;
12'b1100011010110: data = 6'b010101;
12'b1100011010111: data = 6'b010101;
12'b1100011011000: data = 6'b010101;
12'b1100011011001: data = 6'b101010;
12'b1100011011010: data = 6'b101010;
12'b1100011011011: data = 6'b101010;
12'b1100011011100: data = 6'b010101;
12'b1100011011101: data = 6'b000000;
12'b1100011011110: data = 6'b000000;
12'b1100011011111: data = 6'b010101;
12'b1100011100000: data = 6'b010101;
12'b1100011100001: data = 6'b010101;
12'b1100011100010: data = 6'b010101;
12'b1100011100011: data = 6'b010101;
12'b1100011100100: data = 6'b010101;
12'b1100011100101: data = 6'b101001;
12'b1100011100110: data = 6'b101001;
12'b1100011100111: data = 6'b101010;
12'b1100011101000: data = 6'b101010;
12'b1100011101001: data = 6'b101010;
12'b1100011101010: data = 6'b101010;
12'b1100011101011: data = 6'b101010;
12'b1100011101100: data = 6'b101010;
12'b1100011101101: data = 6'b101010;
12'b1100011101110: data = 6'b101010;
12'b1100011101111: data = 6'b101010;
12'b1100011110000: data = 6'b101010;
12'b1100011110001: data = 6'b101010;
12'b1100011110010: data = 6'b101010;
12'b1100011110011: data = 6'b101010;
12'b1100011110100: data = 6'b101010;
12'b1100011110101: data = 6'b111010;
12'b1100011110110: data = 6'b111010;
12'b1100011110111: data = 6'b111110;
12'b1100011111000: data = 6'b111110;
12'b1100011111001: data = 6'b111111;
12'b1100011111010: data = 6'b111111;
12'b1100011111011: data = 6'b111111;
12'b1100011111100: data = 6'b111111;
12'b1100011111101: data = 6'b111111;
12'b1100011111110: data = 6'b111111;
12'b1100011111111: data = 6'b111111;
12'b11000111000000: data = 6'b111111;
12'b11000111000001: data = 6'b111111;
12'b11000111000010: data = 6'b111111;
12'b11000111000011: data = 6'b111111;
12'b11000111000100: data = 6'b111111;
12'b11000111000101: data = 6'b111111;
12'b11000111000110: data = 6'b111111;
12'b11000111000111: data = 6'b111110;
12'b11000111001000: data = 6'b111110;
12'b11000111001001: data = 6'b111110;
12'b11000111001010: data = 6'b111110;
12'b11000111001011: data = 6'b111110;
12'b11000111001100: data = 6'b111010;
12'b11000111001101: data = 6'b111010;
12'b11000111001110: data = 6'b111010;
12'b11000111001111: data = 6'b101010;
12'b11000111010000: data = 6'b101010;
12'b11000111010001: data = 6'b101010;
12'b11000111010010: data = 6'b101010;
12'b11000111010011: data = 6'b101010;
12'b11000111010100: data = 6'b101010;
12'b11000111010101: data = 6'b101010;
12'b11000111010110: data = 6'b101010;
12'b11000111010111: data = 6'b101010;
12'b11000111011000: data = 6'b101010;
12'b11000111011001: data = 6'b101010;
12'b11000111011010: data = 6'b101010;
12'b11000111011011: data = 6'b101010;
12'b11000111011100: data = 6'b101010;
12'b11000111011101: data = 6'b101010;
12'b11000111011110: data = 6'b101010;
12'b11000111011111: data = 6'b101010;
12'b11000111100000: data = 6'b101010;
12'b11000111100001: data = 6'b101010;
12'b11000111100010: data = 6'b101010;
12'b11000111100011: data = 6'b101010;
12'b11000111100100: data = 6'b101010;
12'b11000111100101: data = 6'b101010;
12'b11000111100110: data = 6'b101010;
12'b11000111100111: data = 6'b101010;
12'b11000111101000: data = 6'b101010;
12'b11000111101001: data = 6'b101010;
12'b11000111101010: data = 6'b101010;
12'b11000111101011: data = 6'b101010;
12'b11000111101100: data = 6'b101010;
12'b11000111101101: data = 6'b101010;
12'b11000111101110: data = 6'b101010;
12'b11000111101111: data = 6'b101010;
12'b11000111110000: data = 6'b101010;
12'b11000111110001: data = 6'b101010;
12'b11000111110010: data = 6'b101010;
12'b11000111110011: data = 6'b101010;
12'b11000111110100: data = 6'b101010;
12'b11000111110101: data = 6'b101010;
12'b11000111110110: data = 6'b101010;
12'b11000111110111: data = 6'b101010;
12'b11000111111000: data = 6'b101010;
12'b11000111111001: data = 6'b101001;
12'b11000111111010: data = 6'b101001;
12'b11000111111011: data = 6'b101001;
12'b11000111111100: data = 6'b010101;
12'b11000111111101: data = 6'b010101;
12'b11000111111110: data = 6'b010101;
12'b11000111111111: data = 6'b010101;
12'b110001110000000: data = 6'b010101;
12'b110001110000001: data = 6'b010101;
12'b110001110000010: data = 6'b010101;
12'b110001110000011: data = 6'b010101;
12'b110001110000100: data = 6'b010101;
12'b110001110000101: data = 6'b010101;
12'b110001110000110: data = 6'b010101;
12'b110001110000111: data = 6'b010101;
12'b110001110001000: data = 6'b010101;
12'b110001110001001: data = 6'b010101;
12'b110001110001010: data = 6'b010101;
12'b110001110001011: data = 6'b010101;
12'b110001110001100: data = 6'b000000;
12'b110001110001101: data = 6'b000000;
12'b110001110001110: data = 6'b101010;
12'b110001110001111: data = 6'b101010;
12'b110001110010000: data = 6'b101010;
12'b110001110010001: data = 6'b101010;
12'b110001110010010: data = 6'b010101;
12'b110001110010011: data = 6'b010101;
12'b110001110010100: data = 6'b010101;
12'b110001110010101: data = 6'b010101;
12'b110001110010110: data = 6'b010101;
12'b110001110010111: data = 6'b010101;
12'b110001110011000: data = 6'b010101;
12'b110001110011001: data = 6'b010101;
12'b110001110011010: data = 6'b010101;
12'b110001110011011: data = 6'b010101;
12'b110001110011100: data = 6'b010101;
12'b110001110011101: data = 6'b010101;
12'b110001110011110: data = 6'b010101;
12'b110001110011111: data = 6'b010101;
12'b110001110100000: data = 6'b010101;
12'b110001110100001: data = 6'b010101;
12'b110001110100010: data = 6'b010101;
12'b110001110100011: data = 6'b010101;
12'b110001110100100: data = 6'b010101;
12'b110001110100101: data = 6'b010101;
12'b110001110100110: data = 6'b010101;
12'b110001110100111: data = 6'b010101;
12'b110001110101000: data = 6'b010101;
12'b110001110101001: data = 6'b010101;
12'b110001110101010: data = 6'b010101;
12'b1100100000000: data = 6'b010101;
12'b1100100000001: data = 6'b010101;
12'b1100100000010: data = 6'b010101;
12'b1100100000011: data = 6'b010101;
12'b1100100000100: data = 6'b010101;
12'b1100100000101: data = 6'b010101;
12'b1100100000110: data = 6'b010101;
12'b1100100000111: data = 6'b010101;
12'b1100100001000: data = 6'b010101;
12'b1100100001001: data = 6'b010101;
12'b1100100001010: data = 6'b010101;
12'b1100100001011: data = 6'b010101;
12'b1100100001100: data = 6'b010101;
12'b1100100001101: data = 6'b010101;
12'b1100100001110: data = 6'b010101;
12'b1100100001111: data = 6'b010101;
12'b1100100010000: data = 6'b010101;
12'b1100100010001: data = 6'b010101;
12'b1100100010010: data = 6'b010101;
12'b1100100010011: data = 6'b010101;
12'b1100100010100: data = 6'b010101;
12'b1100100010101: data = 6'b010101;
12'b1100100010110: data = 6'b010101;
12'b1100100010111: data = 6'b010101;
12'b1100100011000: data = 6'b010101;
12'b1100100011001: data = 6'b101010;
12'b1100100011010: data = 6'b101010;
12'b1100100011011: data = 6'b101010;
12'b1100100011100: data = 6'b010101;
12'b1100100011101: data = 6'b000000;
12'b1100100011110: data = 6'b000000;
12'b1100100011111: data = 6'b010101;
12'b1100100100000: data = 6'b010101;
12'b1100100100001: data = 6'b010101;
12'b1100100100010: data = 6'b010101;
12'b1100100100011: data = 6'b010101;
12'b1100100100100: data = 6'b010101;
12'b1100100100101: data = 6'b101001;
12'b1100100100110: data = 6'b101001;
12'b1100100100111: data = 6'b101010;
12'b1100100101000: data = 6'b101010;
12'b1100100101001: data = 6'b101010;
12'b1100100101010: data = 6'b101010;
12'b1100100101011: data = 6'b101010;
12'b1100100101100: data = 6'b101010;
12'b1100100101101: data = 6'b101010;
12'b1100100101110: data = 6'b101010;
12'b1100100101111: data = 6'b101010;
12'b1100100110000: data = 6'b101010;
12'b1100100110001: data = 6'b101010;
12'b1100100110010: data = 6'b101010;
12'b1100100110011: data = 6'b101010;
12'b1100100110100: data = 6'b101010;
12'b1100100110101: data = 6'b111010;
12'b1100100110110: data = 6'b111010;
12'b1100100110111: data = 6'b111110;
12'b1100100111000: data = 6'b111110;
12'b1100100111001: data = 6'b111111;
12'b1100100111010: data = 6'b111111;
12'b1100100111011: data = 6'b111111;
12'b1100100111100: data = 6'b111111;
12'b1100100111101: data = 6'b111111;
12'b1100100111110: data = 6'b111111;
12'b1100100111111: data = 6'b111111;
12'b11001001000000: data = 6'b111111;
12'b11001001000001: data = 6'b111111;
12'b11001001000010: data = 6'b111111;
12'b11001001000011: data = 6'b111111;
12'b11001001000100: data = 6'b111111;
12'b11001001000101: data = 6'b111111;
12'b11001001000110: data = 6'b111111;
12'b11001001000111: data = 6'b111110;
12'b11001001001000: data = 6'b111110;
12'b11001001001001: data = 6'b111110;
12'b11001001001010: data = 6'b111110;
12'b11001001001011: data = 6'b111110;
12'b11001001001100: data = 6'b111010;
12'b11001001001101: data = 6'b111010;
12'b11001001001110: data = 6'b111010;
12'b11001001001111: data = 6'b101010;
12'b11001001010000: data = 6'b101010;
12'b11001001010001: data = 6'b101010;
12'b11001001010010: data = 6'b101010;
12'b11001001010011: data = 6'b101010;
12'b11001001010100: data = 6'b101010;
12'b11001001010101: data = 6'b101010;
12'b11001001010110: data = 6'b101010;
12'b11001001010111: data = 6'b101010;
12'b11001001011000: data = 6'b101010;
12'b11001001011001: data = 6'b101010;
12'b11001001011010: data = 6'b101010;
12'b11001001011011: data = 6'b101010;
12'b11001001011100: data = 6'b101010;
12'b11001001011101: data = 6'b101010;
12'b11001001011110: data = 6'b101010;
12'b11001001011111: data = 6'b101010;
12'b11001001100000: data = 6'b101010;
12'b11001001100001: data = 6'b101010;
12'b11001001100010: data = 6'b101010;
12'b11001001100011: data = 6'b101010;
12'b11001001100100: data = 6'b101010;
12'b11001001100101: data = 6'b101010;
12'b11001001100110: data = 6'b101010;
12'b11001001100111: data = 6'b101010;
12'b11001001101000: data = 6'b101010;
12'b11001001101001: data = 6'b101010;
12'b11001001101010: data = 6'b101010;
12'b11001001101011: data = 6'b101010;
12'b11001001101100: data = 6'b101010;
12'b11001001101101: data = 6'b101010;
12'b11001001101110: data = 6'b101010;
12'b11001001101111: data = 6'b101010;
12'b11001001110000: data = 6'b101010;
12'b11001001110001: data = 6'b101010;
12'b11001001110010: data = 6'b101010;
12'b11001001110011: data = 6'b101010;
12'b11001001110100: data = 6'b101010;
12'b11001001110101: data = 6'b101010;
12'b11001001110110: data = 6'b101010;
12'b11001001110111: data = 6'b101010;
12'b11001001111000: data = 6'b101010;
12'b11001001111001: data = 6'b101001;
12'b11001001111010: data = 6'b101001;
12'b11001001111011: data = 6'b101001;
12'b11001001111100: data = 6'b010101;
12'b11001001111101: data = 6'b101001;
12'b11001001111110: data = 6'b010101;
12'b11001001111111: data = 6'b010101;
12'b110010010000000: data = 6'b010101;
12'b110010010000001: data = 6'b010101;
12'b110010010000010: data = 6'b010101;
12'b110010010000011: data = 6'b010101;
12'b110010010000100: data = 6'b010101;
12'b110010010000101: data = 6'b010101;
12'b110010010000110: data = 6'b010101;
12'b110010010000111: data = 6'b010101;
12'b110010010001000: data = 6'b010101;
12'b110010010001001: data = 6'b010101;
12'b110010010001010: data = 6'b010101;
12'b110010010001011: data = 6'b010101;
12'b110010010001100: data = 6'b000000;
12'b110010010001101: data = 6'b000000;
12'b110010010001110: data = 6'b101010;
12'b110010010001111: data = 6'b101010;
12'b110010010010000: data = 6'b101010;
12'b110010010010001: data = 6'b101010;
12'b110010010010010: data = 6'b010101;
12'b110010010010011: data = 6'b010101;
12'b110010010010100: data = 6'b010101;
12'b110010010010101: data = 6'b010101;
12'b110010010010110: data = 6'b010101;
12'b110010010010111: data = 6'b010101;
12'b110010010011000: data = 6'b010101;
12'b110010010011001: data = 6'b010101;
12'b110010010011010: data = 6'b010101;
12'b110010010011011: data = 6'b010101;
12'b110010010011100: data = 6'b010101;
12'b110010010011101: data = 6'b010101;
12'b110010010011110: data = 6'b010101;
12'b110010010011111: data = 6'b010101;
12'b110010010100000: data = 6'b010101;
12'b110010010100001: data = 6'b010101;
12'b110010010100010: data = 6'b010101;
12'b110010010100011: data = 6'b010101;
12'b110010010100100: data = 6'b010101;
12'b110010010100101: data = 6'b010101;
12'b110010010100110: data = 6'b010101;
12'b110010010100111: data = 6'b010101;
12'b110010010101000: data = 6'b010101;
12'b110010010101001: data = 6'b010101;
12'b110010010101010: data = 6'b010101;
12'b1100101000000: data = 6'b010101;
12'b1100101000001: data = 6'b010101;
12'b1100101000010: data = 6'b010101;
12'b1100101000011: data = 6'b010101;
12'b1100101000100: data = 6'b010101;
12'b1100101000101: data = 6'b010101;
12'b1100101000110: data = 6'b010101;
12'b1100101000111: data = 6'b010101;
12'b1100101001000: data = 6'b010101;
12'b1100101001001: data = 6'b010101;
12'b1100101001010: data = 6'b010101;
12'b1100101001011: data = 6'b010101;
12'b1100101001100: data = 6'b010101;
12'b1100101001101: data = 6'b010101;
12'b1100101001110: data = 6'b010101;
12'b1100101001111: data = 6'b010101;
12'b1100101010000: data = 6'b010101;
12'b1100101010001: data = 6'b010101;
12'b1100101010010: data = 6'b010101;
12'b1100101010011: data = 6'b010101;
12'b1100101010100: data = 6'b010101;
12'b1100101010101: data = 6'b010101;
12'b1100101010110: data = 6'b010101;
12'b1100101010111: data = 6'b010101;
12'b1100101011000: data = 6'b010101;
12'b1100101011001: data = 6'b101010;
12'b1100101011010: data = 6'b101010;
12'b1100101011011: data = 6'b101010;
12'b1100101011100: data = 6'b010101;
12'b1100101011101: data = 6'b000000;
12'b1100101011110: data = 6'b000000;
12'b1100101011111: data = 6'b010101;
12'b1100101100000: data = 6'b010101;
12'b1100101100001: data = 6'b010101;
12'b1100101100010: data = 6'b010101;
12'b1100101100011: data = 6'b010101;
12'b1100101100100: data = 6'b010101;
12'b1100101100101: data = 6'b101001;
12'b1100101100110: data = 6'b101001;
12'b1100101100111: data = 6'b101010;
12'b1100101101000: data = 6'b101010;
12'b1100101101001: data = 6'b101010;
12'b1100101101010: data = 6'b101010;
12'b1100101101011: data = 6'b101010;
12'b1100101101100: data = 6'b101010;
12'b1100101101101: data = 6'b101010;
12'b1100101101110: data = 6'b101010;
12'b1100101101111: data = 6'b101010;
12'b1100101110000: data = 6'b101010;
12'b1100101110001: data = 6'b101010;
12'b1100101110010: data = 6'b101010;
12'b1100101110011: data = 6'b101010;
12'b1100101110100: data = 6'b101010;
12'b1100101110101: data = 6'b111010;
12'b1100101110110: data = 6'b111010;
12'b1100101110111: data = 6'b111110;
12'b1100101111000: data = 6'b111110;
12'b1100101111001: data = 6'b111111;
12'b1100101111010: data = 6'b111111;
12'b1100101111011: data = 6'b111111;
12'b1100101111100: data = 6'b111111;
12'b1100101111101: data = 6'b111111;
12'b1100101111110: data = 6'b111111;
12'b1100101111111: data = 6'b111111;
12'b11001011000000: data = 6'b111111;
12'b11001011000001: data = 6'b111111;
12'b11001011000010: data = 6'b111111;
12'b11001011000011: data = 6'b111111;
12'b11001011000100: data = 6'b111111;
12'b11001011000101: data = 6'b111111;
12'b11001011000110: data = 6'b111111;
12'b11001011000111: data = 6'b111110;
12'b11001011001000: data = 6'b111110;
12'b11001011001001: data = 6'b111110;
12'b11001011001010: data = 6'b111110;
12'b11001011001011: data = 6'b111110;
12'b11001011001100: data = 6'b111010;
12'b11001011001101: data = 6'b111010;
12'b11001011001110: data = 6'b111010;
12'b11001011001111: data = 6'b101010;
12'b11001011010000: data = 6'b101010;
12'b11001011010001: data = 6'b101010;
12'b11001011010010: data = 6'b101010;
12'b11001011010011: data = 6'b101010;
12'b11001011010100: data = 6'b101010;
12'b11001011010101: data = 6'b101010;
12'b11001011010110: data = 6'b101010;
12'b11001011010111: data = 6'b101010;
12'b11001011011000: data = 6'b101010;
12'b11001011011001: data = 6'b101010;
12'b11001011011010: data = 6'b101010;
12'b11001011011011: data = 6'b101010;
12'b11001011011100: data = 6'b101010;
12'b11001011011101: data = 6'b101010;
12'b11001011011110: data = 6'b101010;
12'b11001011011111: data = 6'b101010;
12'b11001011100000: data = 6'b101010;
12'b11001011100001: data = 6'b101010;
12'b11001011100010: data = 6'b101010;
12'b11001011100011: data = 6'b101010;
12'b11001011100100: data = 6'b101010;
12'b11001011100101: data = 6'b101010;
12'b11001011100110: data = 6'b101010;
12'b11001011100111: data = 6'b101010;
12'b11001011101000: data = 6'b101010;
12'b11001011101001: data = 6'b101010;
12'b11001011101010: data = 6'b101010;
12'b11001011101011: data = 6'b101010;
12'b11001011101100: data = 6'b101010;
12'b11001011101101: data = 6'b101010;
12'b11001011101110: data = 6'b101010;
12'b11001011101111: data = 6'b101010;
12'b11001011110000: data = 6'b101010;
12'b11001011110001: data = 6'b101010;
12'b11001011110010: data = 6'b101010;
12'b11001011110011: data = 6'b101010;
12'b11001011110100: data = 6'b101010;
12'b11001011110101: data = 6'b101010;
12'b11001011110110: data = 6'b101010;
12'b11001011110111: data = 6'b101010;
12'b11001011111000: data = 6'b101010;
12'b11001011111001: data = 6'b101001;
12'b11001011111010: data = 6'b101001;
12'b11001011111011: data = 6'b101001;
12'b11001011111100: data = 6'b010101;
12'b11001011111101: data = 6'b010101;
12'b11001011111110: data = 6'b010101;
12'b11001011111111: data = 6'b010101;
12'b110010110000000: data = 6'b010101;
12'b110010110000001: data = 6'b010101;
12'b110010110000010: data = 6'b010101;
12'b110010110000011: data = 6'b010101;
12'b110010110000100: data = 6'b010101;
12'b110010110000101: data = 6'b010101;
12'b110010110000110: data = 6'b010101;
12'b110010110000111: data = 6'b010101;
12'b110010110001000: data = 6'b010101;
12'b110010110001001: data = 6'b010101;
12'b110010110001010: data = 6'b010101;
12'b110010110001011: data = 6'b010101;
12'b110010110001100: data = 6'b000000;
12'b110010110001101: data = 6'b000000;
12'b110010110001110: data = 6'b101010;
12'b110010110001111: data = 6'b101010;
12'b110010110010000: data = 6'b101010;
12'b110010110010001: data = 6'b101010;
12'b110010110010010: data = 6'b010101;
12'b110010110010011: data = 6'b010101;
12'b110010110010100: data = 6'b010101;
12'b110010110010101: data = 6'b010101;
12'b110010110010110: data = 6'b010101;
12'b110010110010111: data = 6'b010101;
12'b110010110011000: data = 6'b010101;
12'b110010110011001: data = 6'b010101;
12'b110010110011010: data = 6'b010101;
12'b110010110011011: data = 6'b010101;
12'b110010110011100: data = 6'b010101;
12'b110010110011101: data = 6'b010101;
12'b110010110011110: data = 6'b010101;
12'b110010110011111: data = 6'b010101;
12'b110010110100000: data = 6'b010101;
12'b110010110100001: data = 6'b010101;
12'b110010110100010: data = 6'b010101;
12'b110010110100011: data = 6'b010101;
12'b110010110100100: data = 6'b010101;
12'b110010110100101: data = 6'b010101;
12'b110010110100110: data = 6'b010101;
12'b110010110100111: data = 6'b010101;
12'b110010110101000: data = 6'b010101;
12'b110010110101001: data = 6'b010101;
12'b110010110101010: data = 6'b010101;
12'b1100110000000: data = 6'b010101;
12'b1100110000001: data = 6'b010101;
12'b1100110000010: data = 6'b010101;
12'b1100110000011: data = 6'b010101;
12'b1100110000100: data = 6'b010101;
12'b1100110000101: data = 6'b010101;
12'b1100110000110: data = 6'b010101;
12'b1100110000111: data = 6'b010101;
12'b1100110001000: data = 6'b010101;
12'b1100110001001: data = 6'b010101;
12'b1100110001010: data = 6'b010101;
12'b1100110001011: data = 6'b010101;
12'b1100110001100: data = 6'b010101;
12'b1100110001101: data = 6'b010101;
12'b1100110001110: data = 6'b010101;
12'b1100110001111: data = 6'b010101;
12'b1100110010000: data = 6'b010101;
12'b1100110010001: data = 6'b010101;
12'b1100110010010: data = 6'b010101;
12'b1100110010011: data = 6'b010101;
12'b1100110010100: data = 6'b010101;
12'b1100110010101: data = 6'b010101;
12'b1100110010110: data = 6'b010101;
12'b1100110010111: data = 6'b010101;
12'b1100110011000: data = 6'b010101;
12'b1100110011001: data = 6'b101010;
12'b1100110011010: data = 6'b101010;
12'b1100110011011: data = 6'b101010;
12'b1100110011100: data = 6'b010101;
12'b1100110011101: data = 6'b000000;
12'b1100110011110: data = 6'b000000;
12'b1100110011111: data = 6'b010101;
12'b1100110100000: data = 6'b010101;
12'b1100110100001: data = 6'b010101;
12'b1100110100010: data = 6'b010101;
12'b1100110100011: data = 6'b010101;
12'b1100110100100: data = 6'b010101;
12'b1100110100101: data = 6'b101001;
12'b1100110100110: data = 6'b101001;
12'b1100110100111: data = 6'b101010;
12'b1100110101000: data = 6'b101010;
12'b1100110101001: data = 6'b101010;
12'b1100110101010: data = 6'b101010;
12'b1100110101011: data = 6'b101010;
12'b1100110101100: data = 6'b101010;
12'b1100110101101: data = 6'b101010;
12'b1100110101110: data = 6'b101010;
12'b1100110101111: data = 6'b101010;
12'b1100110110000: data = 6'b101010;
12'b1100110110001: data = 6'b101010;
12'b1100110110010: data = 6'b101010;
12'b1100110110011: data = 6'b101010;
12'b1100110110100: data = 6'b101010;
12'b1100110110101: data = 6'b111010;
12'b1100110110110: data = 6'b111010;
12'b1100110110111: data = 6'b111110;
12'b1100110111000: data = 6'b111111;
12'b1100110111001: data = 6'b111111;
12'b1100110111010: data = 6'b111111;
12'b1100110111011: data = 6'b111111;
12'b1100110111100: data = 6'b111111;
12'b1100110111101: data = 6'b111111;
12'b1100110111110: data = 6'b111111;
12'b1100110111111: data = 6'b111111;
12'b11001101000000: data = 6'b111111;
12'b11001101000001: data = 6'b111111;
12'b11001101000010: data = 6'b111111;
12'b11001101000011: data = 6'b111111;
12'b11001101000100: data = 6'b111111;
12'b11001101000101: data = 6'b111111;
12'b11001101000110: data = 6'b111111;
12'b11001101000111: data = 6'b111111;
12'b11001101001000: data = 6'b111111;
12'b11001101001001: data = 6'b111110;
12'b11001101001010: data = 6'b111110;
12'b11001101001011: data = 6'b111110;
12'b11001101001100: data = 6'b111010;
12'b11001101001101: data = 6'b111010;
12'b11001101001110: data = 6'b111010;
12'b11001101001111: data = 6'b101010;
12'b11001101010000: data = 6'b101010;
12'b11001101010001: data = 6'b101010;
12'b11001101010010: data = 6'b101010;
12'b11001101010011: data = 6'b101010;
12'b11001101010100: data = 6'b101010;
12'b11001101010101: data = 6'b101010;
12'b11001101010110: data = 6'b101010;
12'b11001101010111: data = 6'b101010;
12'b11001101011000: data = 6'b101010;
12'b11001101011001: data = 6'b101010;
12'b11001101011010: data = 6'b101010;
12'b11001101011011: data = 6'b101010;
12'b11001101011100: data = 6'b101010;
12'b11001101011101: data = 6'b101010;
12'b11001101011110: data = 6'b101010;
12'b11001101011111: data = 6'b101010;
12'b11001101100000: data = 6'b101010;
12'b11001101100001: data = 6'b101010;
12'b11001101100010: data = 6'b101010;
12'b11001101100011: data = 6'b101010;
12'b11001101100100: data = 6'b101010;
12'b11001101100101: data = 6'b101010;
12'b11001101100110: data = 6'b101010;
12'b11001101100111: data = 6'b101010;
12'b11001101101000: data = 6'b101010;
12'b11001101101001: data = 6'b101010;
12'b11001101101010: data = 6'b101010;
12'b11001101101011: data = 6'b101010;
12'b11001101101100: data = 6'b101010;
12'b11001101101101: data = 6'b101010;
12'b11001101101110: data = 6'b101010;
12'b11001101101111: data = 6'b101010;
12'b11001101110000: data = 6'b101010;
12'b11001101110001: data = 6'b101010;
12'b11001101110010: data = 6'b101010;
12'b11001101110011: data = 6'b101010;
12'b11001101110100: data = 6'b101010;
12'b11001101110101: data = 6'b101010;
12'b11001101110110: data = 6'b101010;
12'b11001101110111: data = 6'b101010;
12'b11001101111000: data = 6'b101010;
12'b11001101111001: data = 6'b101001;
12'b11001101111010: data = 6'b101001;
12'b11001101111011: data = 6'b101001;
12'b11001101111100: data = 6'b010101;
12'b11001101111101: data = 6'b010101;
12'b11001101111110: data = 6'b010101;
12'b11001101111111: data = 6'b010101;
12'b110011010000000: data = 6'b010101;
12'b110011010000001: data = 6'b010101;
12'b110011010000010: data = 6'b010101;
12'b110011010000011: data = 6'b010101;
12'b110011010000100: data = 6'b010101;
12'b110011010000101: data = 6'b010101;
12'b110011010000110: data = 6'b010101;
12'b110011010000111: data = 6'b010101;
12'b110011010001000: data = 6'b010101;
12'b110011010001001: data = 6'b010101;
12'b110011010001010: data = 6'b010101;
12'b110011010001011: data = 6'b010101;
12'b110011010001100: data = 6'b000000;
12'b110011010001101: data = 6'b000000;
12'b110011010001110: data = 6'b101010;
12'b110011010001111: data = 6'b101010;
12'b110011010010000: data = 6'b101010;
12'b110011010010001: data = 6'b101010;
12'b110011010010010: data = 6'b010101;
12'b110011010010011: data = 6'b010101;
12'b110011010010100: data = 6'b010101;
12'b110011010010101: data = 6'b010101;
12'b110011010010110: data = 6'b010101;
12'b110011010010111: data = 6'b010101;
12'b110011010011000: data = 6'b010101;
12'b110011010011001: data = 6'b010101;
12'b110011010011010: data = 6'b010101;
12'b110011010011011: data = 6'b010101;
12'b110011010011100: data = 6'b010101;
12'b110011010011101: data = 6'b010101;
12'b110011010011110: data = 6'b010101;
12'b110011010011111: data = 6'b010101;
12'b110011010100000: data = 6'b010101;
12'b110011010100001: data = 6'b010101;
12'b110011010100010: data = 6'b010101;
12'b110011010100011: data = 6'b010101;
12'b110011010100100: data = 6'b010101;
12'b110011010100101: data = 6'b010101;
12'b110011010100110: data = 6'b010101;
12'b110011010100111: data = 6'b010101;
12'b110011010101000: data = 6'b010101;
12'b110011010101001: data = 6'b010101;
12'b110011010101010: data = 6'b010101;
12'b1100111000000: data = 6'b010101;
12'b1100111000001: data = 6'b010101;
12'b1100111000010: data = 6'b010101;
12'b1100111000011: data = 6'b010101;
12'b1100111000100: data = 6'b010101;
12'b1100111000101: data = 6'b010101;
12'b1100111000110: data = 6'b010101;
12'b1100111000111: data = 6'b010101;
12'b1100111001000: data = 6'b010101;
12'b1100111001001: data = 6'b010101;
12'b1100111001010: data = 6'b010101;
12'b1100111001011: data = 6'b010101;
12'b1100111001100: data = 6'b010101;
12'b1100111001101: data = 6'b010101;
12'b1100111001110: data = 6'b010101;
12'b1100111001111: data = 6'b010101;
12'b1100111010000: data = 6'b010101;
12'b1100111010001: data = 6'b010101;
12'b1100111010010: data = 6'b010101;
12'b1100111010011: data = 6'b010101;
12'b1100111010100: data = 6'b010101;
12'b1100111010101: data = 6'b010101;
12'b1100111010110: data = 6'b010101;
12'b1100111010111: data = 6'b010101;
12'b1100111011000: data = 6'b010101;
12'b1100111011001: data = 6'b101010;
12'b1100111011010: data = 6'b101010;
12'b1100111011011: data = 6'b101010;
12'b1100111011100: data = 6'b010101;
12'b1100111011101: data = 6'b000000;
12'b1100111011110: data = 6'b000000;
12'b1100111011111: data = 6'b010101;
12'b1100111100000: data = 6'b010101;
12'b1100111100001: data = 6'b010101;
12'b1100111100010: data = 6'b010101;
12'b1100111100011: data = 6'b010101;
12'b1100111100100: data = 6'b010101;
12'b1100111100101: data = 6'b010101;
12'b1100111100110: data = 6'b010101;
12'b1100111100111: data = 6'b010101;
12'b1100111101000: data = 6'b010101;
12'b1100111101001: data = 6'b010101;
12'b1100111101010: data = 6'b101001;
12'b1100111101011: data = 6'b101010;
12'b1100111101100: data = 6'b101010;
12'b1100111101101: data = 6'b101010;
12'b1100111101110: data = 6'b101010;
12'b1100111101111: data = 6'b101010;
12'b1100111110000: data = 6'b101010;
12'b1100111110001: data = 6'b101010;
12'b1100111110010: data = 6'b101010;
12'b1100111110011: data = 6'b101010;
12'b1100111110100: data = 6'b101010;
12'b1100111110101: data = 6'b101010;
12'b1100111110110: data = 6'b101010;
12'b1100111110111: data = 6'b101010;
12'b1100111111000: data = 6'b101010;
12'b1100111111001: data = 6'b101010;
12'b1100111111010: data = 6'b101010;
12'b1100111111011: data = 6'b101010;
12'b1100111111100: data = 6'b101010;
12'b1100111111101: data = 6'b111010;
12'b1100111111110: data = 6'b101010;
12'b1100111111111: data = 6'b101010;
12'b11001111000000: data = 6'b101010;
12'b11001111000001: data = 6'b101010;
12'b11001111000010: data = 6'b101010;
12'b11001111000011: data = 6'b101010;
12'b11001111000100: data = 6'b101010;
12'b11001111000101: data = 6'b101010;
12'b11001111000110: data = 6'b101010;
12'b11001111000111: data = 6'b101010;
12'b11001111001000: data = 6'b101010;
12'b11001111001001: data = 6'b101010;
12'b11001111001010: data = 6'b101010;
12'b11001111001011: data = 6'b101010;
12'b11001111001100: data = 6'b101010;
12'b11001111001101: data = 6'b101010;
12'b11001111001110: data = 6'b101010;
12'b11001111001111: data = 6'b101010;
12'b11001111010000: data = 6'b101010;
12'b11001111010001: data = 6'b101010;
12'b11001111010010: data = 6'b101010;
12'b11001111010011: data = 6'b101010;
12'b11001111010100: data = 6'b101010;
12'b11001111010101: data = 6'b101010;
12'b11001111010110: data = 6'b101010;
12'b11001111010111: data = 6'b101010;
12'b11001111011000: data = 6'b101010;
12'b11001111011001: data = 6'b101010;
12'b11001111011010: data = 6'b101010;
12'b11001111011011: data = 6'b101010;
12'b11001111011100: data = 6'b101010;
12'b11001111011101: data = 6'b101010;
12'b11001111011110: data = 6'b101010;
12'b11001111011111: data = 6'b101010;
12'b11001111100000: data = 6'b101010;
12'b11001111100001: data = 6'b101010;
12'b11001111100010: data = 6'b101010;
12'b11001111100011: data = 6'b101010;
12'b11001111100100: data = 6'b101010;
12'b11001111100101: data = 6'b101010;
12'b11001111100110: data = 6'b101010;
12'b11001111100111: data = 6'b101010;
12'b11001111101000: data = 6'b101010;
12'b11001111101001: data = 6'b101010;
12'b11001111101010: data = 6'b101010;
12'b11001111101011: data = 6'b101010;
12'b11001111101100: data = 6'b101001;
12'b11001111101101: data = 6'b101001;
12'b11001111101110: data = 6'b101001;
12'b11001111101111: data = 6'b101001;
12'b11001111110000: data = 6'b101001;
12'b11001111110001: data = 6'b010101;
12'b11001111110010: data = 6'b010101;
12'b11001111110011: data = 6'b010101;
12'b11001111110100: data = 6'b010101;
12'b11001111110101: data = 6'b010101;
12'b11001111110110: data = 6'b010101;
12'b11001111110111: data = 6'b010101;
12'b11001111111000: data = 6'b010101;
12'b11001111111001: data = 6'b010101;
12'b11001111111010: data = 6'b010101;
12'b11001111111011: data = 6'b010101;
12'b11001111111100: data = 6'b010101;
12'b11001111111101: data = 6'b010101;
12'b11001111111110: data = 6'b010101;
12'b11001111111111: data = 6'b010101;
12'b110011110000000: data = 6'b010101;
12'b110011110000001: data = 6'b010101;
12'b110011110000010: data = 6'b010101;
12'b110011110000011: data = 6'b010101;
12'b110011110000100: data = 6'b010101;
12'b110011110000101: data = 6'b010101;
12'b110011110000110: data = 6'b010101;
12'b110011110000111: data = 6'b010101;
12'b110011110001000: data = 6'b010101;
12'b110011110001001: data = 6'b010101;
12'b110011110001010: data = 6'b010101;
12'b110011110001011: data = 6'b010101;
12'b110011110001100: data = 6'b000000;
12'b110011110001101: data = 6'b000000;
12'b110011110001110: data = 6'b101010;
12'b110011110001111: data = 6'b101010;
12'b110011110010000: data = 6'b101010;
12'b110011110010001: data = 6'b101010;
12'b110011110010010: data = 6'b010101;
12'b110011110010011: data = 6'b010101;
12'b110011110010100: data = 6'b010101;
12'b110011110010101: data = 6'b010101;
12'b110011110010110: data = 6'b010101;
12'b110011110010111: data = 6'b010101;
12'b110011110011000: data = 6'b010101;
12'b110011110011001: data = 6'b010101;
12'b110011110011010: data = 6'b010101;
12'b110011110011011: data = 6'b010101;
12'b110011110011100: data = 6'b010101;
12'b110011110011101: data = 6'b010101;
12'b110011110011110: data = 6'b010101;
12'b110011110011111: data = 6'b010101;
12'b110011110100000: data = 6'b010101;
12'b110011110100001: data = 6'b010101;
12'b110011110100010: data = 6'b010101;
12'b110011110100011: data = 6'b010101;
12'b110011110100100: data = 6'b010101;
12'b110011110100101: data = 6'b010101;
12'b110011110100110: data = 6'b010101;
12'b110011110100111: data = 6'b010101;
12'b110011110101000: data = 6'b010101;
12'b110011110101001: data = 6'b010101;
12'b110011110101010: data = 6'b010101;
12'b1101000000000: data = 6'b010101;
12'b1101000000001: data = 6'b010101;
12'b1101000000010: data = 6'b010101;
12'b1101000000011: data = 6'b010101;
12'b1101000000100: data = 6'b010101;
12'b1101000000101: data = 6'b010101;
12'b1101000000110: data = 6'b010101;
12'b1101000000111: data = 6'b010101;
12'b1101000001000: data = 6'b010101;
12'b1101000001001: data = 6'b010101;
12'b1101000001010: data = 6'b010101;
12'b1101000001011: data = 6'b010101;
12'b1101000001100: data = 6'b010101;
12'b1101000001101: data = 6'b010101;
12'b1101000001110: data = 6'b010101;
12'b1101000001111: data = 6'b010101;
12'b1101000010000: data = 6'b010101;
12'b1101000010001: data = 6'b010101;
12'b1101000010010: data = 6'b010101;
12'b1101000010011: data = 6'b010101;
12'b1101000010100: data = 6'b010101;
12'b1101000010101: data = 6'b010101;
12'b1101000010110: data = 6'b010101;
12'b1101000010111: data = 6'b010101;
12'b1101000011000: data = 6'b010101;
12'b1101000011001: data = 6'b101010;
12'b1101000011010: data = 6'b101010;
12'b1101000011011: data = 6'b101010;
12'b1101000011100: data = 6'b010101;
12'b1101000011101: data = 6'b000000;
12'b1101000011110: data = 6'b000000;
12'b1101000011111: data = 6'b010101;
12'b1101000100000: data = 6'b010101;
12'b1101000100001: data = 6'b010101;
12'b1101000100010: data = 6'b010101;
12'b1101000100011: data = 6'b010101;
12'b1101000100100: data = 6'b010101;
12'b1101000100101: data = 6'b010101;
12'b1101000100110: data = 6'b010101;
12'b1101000100111: data = 6'b000000;
12'b1101000101000: data = 6'b000000;
12'b1101000101001: data = 6'b000000;
12'b1101000101010: data = 6'b000000;
12'b1101000101011: data = 6'b000000;
12'b1101000101100: data = 6'b000000;
12'b1101000101101: data = 6'b000000;
12'b1101000101110: data = 6'b000000;
12'b1101000101111: data = 6'b000000;
12'b1101000110000: data = 6'b000000;
12'b1101000110001: data = 6'b000000;
12'b1101000110010: data = 6'b000000;
12'b1101000110011: data = 6'b000000;
12'b1101000110100: data = 6'b000000;
12'b1101000110101: data = 6'b000000;
12'b1101000110110: data = 6'b000000;
12'b1101000110111: data = 6'b000000;
12'b1101000111000: data = 6'b000000;
12'b1101000111001: data = 6'b000000;
12'b1101000111010: data = 6'b000000;
12'b1101000111011: data = 6'b000000;
12'b1101000111100: data = 6'b000000;
12'b1101000111101: data = 6'b000000;
12'b1101000111110: data = 6'b000000;
12'b1101000111111: data = 6'b000000;
12'b11010001000000: data = 6'b000000;
12'b11010001000001: data = 6'b000000;
12'b11010001000010: data = 6'b000000;
12'b11010001000011: data = 6'b000000;
12'b11010001000100: data = 6'b000000;
12'b11010001000101: data = 6'b000000;
12'b11010001000110: data = 6'b000000;
12'b11010001000111: data = 6'b000000;
12'b11010001001000: data = 6'b000000;
12'b11010001001001: data = 6'b000000;
12'b11010001001010: data = 6'b000000;
12'b11010001001011: data = 6'b000000;
12'b11010001001100: data = 6'b000000;
12'b11010001001101: data = 6'b000000;
12'b11010001001110: data = 6'b000000;
12'b11010001001111: data = 6'b000000;
12'b11010001010000: data = 6'b000000;
12'b11010001010001: data = 6'b000000;
12'b11010001010010: data = 6'b000000;
12'b11010001010011: data = 6'b000000;
12'b11010001010100: data = 6'b000000;
12'b11010001010101: data = 6'b000000;
12'b11010001010110: data = 6'b000000;
12'b11010001010111: data = 6'b000000;
12'b11010001011000: data = 6'b000000;
12'b11010001011001: data = 6'b000000;
12'b11010001011010: data = 6'b000000;
12'b11010001011011: data = 6'b000000;
12'b11010001011100: data = 6'b000000;
12'b11010001011101: data = 6'b000000;
12'b11010001011110: data = 6'b000000;
12'b11010001011111: data = 6'b000000;
12'b11010001100000: data = 6'b000000;
12'b11010001100001: data = 6'b000000;
12'b11010001100010: data = 6'b000000;
12'b11010001100011: data = 6'b000000;
12'b11010001100100: data = 6'b000000;
12'b11010001100101: data = 6'b000000;
12'b11010001100110: data = 6'b000000;
12'b11010001100111: data = 6'b000000;
12'b11010001101000: data = 6'b000000;
12'b11010001101001: data = 6'b000000;
12'b11010001101010: data = 6'b000000;
12'b11010001101011: data = 6'b000000;
12'b11010001101100: data = 6'b000000;
12'b11010001101101: data = 6'b000000;
12'b11010001101110: data = 6'b000000;
12'b11010001101111: data = 6'b000000;
12'b11010001110000: data = 6'b000000;
12'b11010001110001: data = 6'b000000;
12'b11010001110010: data = 6'b000000;
12'b11010001110011: data = 6'b000000;
12'b11010001110100: data = 6'b000000;
12'b11010001110101: data = 6'b000000;
12'b11010001110110: data = 6'b000000;
12'b11010001110111: data = 6'b000000;
12'b11010001111000: data = 6'b000000;
12'b11010001111001: data = 6'b000000;
12'b11010001111010: data = 6'b000000;
12'b11010001111011: data = 6'b000000;
12'b11010001111100: data = 6'b000000;
12'b11010001111101: data = 6'b000000;
12'b11010001111110: data = 6'b000000;
12'b11010001111111: data = 6'b000000;
12'b110100010000000: data = 6'b000000;
12'b110100010000001: data = 6'b000000;
12'b110100010000010: data = 6'b000000;
12'b110100010000011: data = 6'b000000;
12'b110100010000100: data = 6'b010101;
12'b110100010000101: data = 6'b010101;
12'b110100010000110: data = 6'b010101;
12'b110100010000111: data = 6'b010101;
12'b110100010001000: data = 6'b010101;
12'b110100010001001: data = 6'b010101;
12'b110100010001010: data = 6'b010101;
12'b110100010001011: data = 6'b010101;
12'b110100010001100: data = 6'b000000;
12'b110100010001101: data = 6'b000000;
12'b110100010001110: data = 6'b101010;
12'b110100010001111: data = 6'b101010;
12'b110100010010000: data = 6'b101010;
12'b110100010010001: data = 6'b101010;
12'b110100010010010: data = 6'b010101;
12'b110100010010011: data = 6'b010101;
12'b110100010010100: data = 6'b010101;
12'b110100010010101: data = 6'b010101;
12'b110100010010110: data = 6'b010101;
12'b110100010010111: data = 6'b010101;
12'b110100010011000: data = 6'b010101;
12'b110100010011001: data = 6'b010101;
12'b110100010011010: data = 6'b010101;
12'b110100010011011: data = 6'b010101;
12'b110100010011100: data = 6'b010101;
12'b110100010011101: data = 6'b010101;
12'b110100010011110: data = 6'b010101;
12'b110100010011111: data = 6'b010101;
12'b110100010100000: data = 6'b010101;
12'b110100010100001: data = 6'b010101;
12'b110100010100010: data = 6'b010101;
12'b110100010100011: data = 6'b010101;
12'b110100010100100: data = 6'b010101;
12'b110100010100101: data = 6'b010101;
12'b110100010100110: data = 6'b010101;
12'b110100010100111: data = 6'b010101;
12'b110100010101000: data = 6'b010101;
12'b110100010101001: data = 6'b010101;
12'b110100010101010: data = 6'b010101;
12'b1101001000000: data = 6'b010101;
12'b1101001000001: data = 6'b010101;
12'b1101001000010: data = 6'b010101;
12'b1101001000011: data = 6'b010101;
12'b1101001000100: data = 6'b010101;
12'b1101001000101: data = 6'b010101;
12'b1101001000110: data = 6'b010101;
12'b1101001000111: data = 6'b010101;
12'b1101001001000: data = 6'b010101;
12'b1101001001001: data = 6'b010101;
12'b1101001001010: data = 6'b010101;
12'b1101001001011: data = 6'b010101;
12'b1101001001100: data = 6'b010101;
12'b1101001001101: data = 6'b010101;
12'b1101001001110: data = 6'b010101;
12'b1101001001111: data = 6'b010101;
12'b1101001010000: data = 6'b010101;
12'b1101001010001: data = 6'b010101;
12'b1101001010010: data = 6'b010101;
12'b1101001010011: data = 6'b010101;
12'b1101001010100: data = 6'b010101;
12'b1101001010101: data = 6'b010101;
12'b1101001010110: data = 6'b010101;
12'b1101001010111: data = 6'b010101;
12'b1101001011000: data = 6'b010101;
12'b1101001011001: data = 6'b101010;
12'b1101001011010: data = 6'b101010;
12'b1101001011011: data = 6'b101010;
12'b1101001011100: data = 6'b010101;
12'b1101001011101: data = 6'b000000;
12'b1101001011110: data = 6'b000000;
12'b1101001011111: data = 6'b010101;
12'b1101001100000: data = 6'b010101;
12'b1101001100001: data = 6'b010101;
12'b1101001100010: data = 6'b010101;
12'b1101001100011: data = 6'b010101;
12'b1101001100100: data = 6'b010101;
12'b1101001100101: data = 6'b010101;
12'b1101001100110: data = 6'b010101;
12'b1101001100111: data = 6'b000000;
12'b1101001101000: data = 6'b000000;
12'b1101001101001: data = 6'b000000;
12'b1101001101010: data = 6'b000000;
12'b1101001101011: data = 6'b000000;
12'b1101001101100: data = 6'b000000;
12'b1101001101101: data = 6'b000000;
12'b1101001101110: data = 6'b000000;
12'b1101001101111: data = 6'b000000;
12'b1101001110000: data = 6'b000000;
12'b1101001110001: data = 6'b000000;
12'b1101001110010: data = 6'b000000;
12'b1101001110011: data = 6'b000000;
12'b1101001110100: data = 6'b000000;
12'b1101001110101: data = 6'b000000;
12'b1101001110110: data = 6'b000000;
12'b1101001110111: data = 6'b000000;
12'b1101001111000: data = 6'b000000;
12'b1101001111001: data = 6'b000000;
12'b1101001111010: data = 6'b000000;
12'b1101001111011: data = 6'b000000;
12'b1101001111100: data = 6'b000000;
12'b1101001111101: data = 6'b000000;
12'b1101001111110: data = 6'b000000;
12'b1101001111111: data = 6'b000000;
12'b11010011000000: data = 6'b000000;
12'b11010011000001: data = 6'b000000;
12'b11010011000010: data = 6'b000000;
12'b11010011000011: data = 6'b000000;
12'b11010011000100: data = 6'b000000;
12'b11010011000101: data = 6'b000000;
12'b11010011000110: data = 6'b000000;
12'b11010011000111: data = 6'b000000;
12'b11010011001000: data = 6'b000000;
12'b11010011001001: data = 6'b000000;
12'b11010011001010: data = 6'b000000;
12'b11010011001011: data = 6'b000000;
12'b11010011001100: data = 6'b000000;
12'b11010011001101: data = 6'b000000;
12'b11010011001110: data = 6'b000000;
12'b11010011001111: data = 6'b000000;
12'b11010011010000: data = 6'b000000;
12'b11010011010001: data = 6'b000000;
12'b11010011010010: data = 6'b000000;
12'b11010011010011: data = 6'b000000;
12'b11010011010100: data = 6'b000000;
12'b11010011010101: data = 6'b000000;
12'b11010011010110: data = 6'b000000;
12'b11010011010111: data = 6'b000000;
12'b11010011011000: data = 6'b000000;
12'b11010011011001: data = 6'b000000;
12'b11010011011010: data = 6'b000000;
12'b11010011011011: data = 6'b000000;
12'b11010011011100: data = 6'b000000;
12'b11010011011101: data = 6'b000000;
12'b11010011011110: data = 6'b000000;
12'b11010011011111: data = 6'b000000;
12'b11010011100000: data = 6'b000000;
12'b11010011100001: data = 6'b000000;
12'b11010011100010: data = 6'b000000;
12'b11010011100011: data = 6'b000000;
12'b11010011100100: data = 6'b000000;
12'b11010011100101: data = 6'b000000;
12'b11010011100110: data = 6'b000000;
12'b11010011100111: data = 6'b000000;
12'b11010011101000: data = 6'b000000;
12'b11010011101001: data = 6'b000000;
12'b11010011101010: data = 6'b000000;
12'b11010011101011: data = 6'b000000;
12'b11010011101100: data = 6'b000000;
12'b11010011101101: data = 6'b000000;
12'b11010011101110: data = 6'b000000;
12'b11010011101111: data = 6'b000000;
12'b11010011110000: data = 6'b000000;
12'b11010011110001: data = 6'b000000;
12'b11010011110010: data = 6'b000000;
12'b11010011110011: data = 6'b000000;
12'b11010011110100: data = 6'b000000;
12'b11010011110101: data = 6'b000000;
12'b11010011110110: data = 6'b000000;
12'b11010011110111: data = 6'b000000;
12'b11010011111000: data = 6'b000000;
12'b11010011111001: data = 6'b000000;
12'b11010011111010: data = 6'b000000;
12'b11010011111011: data = 6'b000000;
12'b11010011111100: data = 6'b000000;
12'b11010011111101: data = 6'b000000;
12'b11010011111110: data = 6'b000000;
12'b11010011111111: data = 6'b000000;
12'b110100110000000: data = 6'b000000;
12'b110100110000001: data = 6'b000000;
12'b110100110000010: data = 6'b000000;
12'b110100110000011: data = 6'b000000;
12'b110100110000100: data = 6'b010101;
12'b110100110000101: data = 6'b010101;
12'b110100110000110: data = 6'b010101;
12'b110100110000111: data = 6'b010101;
12'b110100110001000: data = 6'b010101;
12'b110100110001001: data = 6'b010101;
12'b110100110001010: data = 6'b010101;
12'b110100110001011: data = 6'b010101;
12'b110100110001100: data = 6'b000000;
12'b110100110001101: data = 6'b000000;
12'b110100110001110: data = 6'b101010;
12'b110100110001111: data = 6'b101010;
12'b110100110010000: data = 6'b101010;
12'b110100110010001: data = 6'b101010;
12'b110100110010010: data = 6'b010101;
12'b110100110010011: data = 6'b010101;
12'b110100110010100: data = 6'b010101;
12'b110100110010101: data = 6'b010101;
12'b110100110010110: data = 6'b010101;
12'b110100110010111: data = 6'b010101;
12'b110100110011000: data = 6'b010101;
12'b110100110011001: data = 6'b010101;
12'b110100110011010: data = 6'b010101;
12'b110100110011011: data = 6'b010101;
12'b110100110011100: data = 6'b010101;
12'b110100110011101: data = 6'b010101;
12'b110100110011110: data = 6'b010101;
12'b110100110011111: data = 6'b010101;
12'b110100110100000: data = 6'b010101;
12'b110100110100001: data = 6'b010101;
12'b110100110100010: data = 6'b010101;
12'b110100110100011: data = 6'b010101;
12'b110100110100100: data = 6'b010101;
12'b110100110100101: data = 6'b010101;
12'b110100110100110: data = 6'b010101;
12'b110100110100111: data = 6'b010101;
12'b110100110101000: data = 6'b010101;
12'b110100110101001: data = 6'b010101;
12'b110100110101010: data = 6'b010101;
12'b1101010000000: data = 6'b010101;
12'b1101010000001: data = 6'b010101;
12'b1101010000010: data = 6'b010101;
12'b1101010000011: data = 6'b010101;
12'b1101010000100: data = 6'b010101;
12'b1101010000101: data = 6'b010101;
12'b1101010000110: data = 6'b010101;
12'b1101010000111: data = 6'b010101;
12'b1101010001000: data = 6'b010101;
12'b1101010001001: data = 6'b010101;
12'b1101010001010: data = 6'b010101;
12'b1101010001011: data = 6'b010101;
12'b1101010001100: data = 6'b010101;
12'b1101010001101: data = 6'b010101;
12'b1101010001110: data = 6'b010101;
12'b1101010001111: data = 6'b010101;
12'b1101010010000: data = 6'b010101;
12'b1101010010001: data = 6'b010101;
12'b1101010010010: data = 6'b010101;
12'b1101010010011: data = 6'b010101;
12'b1101010010100: data = 6'b010101;
12'b1101010010101: data = 6'b010101;
12'b1101010010110: data = 6'b010101;
12'b1101010010111: data = 6'b010101;
12'b1101010011000: data = 6'b010101;
12'b1101010011001: data = 6'b101010;
12'b1101010011010: data = 6'b101010;
12'b1101010011011: data = 6'b101010;
12'b1101010011100: data = 6'b101010;
12'b1101010011101: data = 6'b010101;
12'b1101010011110: data = 6'b010101;
12'b1101010011111: data = 6'b010101;
12'b1101010100000: data = 6'b010101;
12'b1101010100001: data = 6'b010101;
12'b1101010100010: data = 6'b010101;
12'b1101010100011: data = 6'b010101;
12'b1101010100100: data = 6'b010101;
12'b1101010100101: data = 6'b010101;
12'b1101010100110: data = 6'b010101;
12'b1101010100111: data = 6'b000000;
12'b1101010101000: data = 6'b000000;
12'b1101010101001: data = 6'b000000;
12'b1101010101010: data = 6'b000000;
12'b1101010101011: data = 6'b000000;
12'b1101010101100: data = 6'b000000;
12'b1101010101101: data = 6'b000000;
12'b1101010101110: data = 6'b000000;
12'b1101010101111: data = 6'b000000;
12'b1101010110000: data = 6'b000000;
12'b1101010110001: data = 6'b000000;
12'b1101010110010: data = 6'b000000;
12'b1101010110011: data = 6'b000000;
12'b1101010110100: data = 6'b000000;
12'b1101010110101: data = 6'b000000;
12'b1101010110110: data = 6'b000000;
12'b1101010110111: data = 6'b000000;
12'b1101010111000: data = 6'b000000;
12'b1101010111001: data = 6'b000000;
12'b1101010111010: data = 6'b000000;
12'b1101010111011: data = 6'b000000;
12'b1101010111100: data = 6'b000000;
12'b1101010111101: data = 6'b000000;
12'b1101010111110: data = 6'b000000;
12'b1101010111111: data = 6'b000000;
12'b11010101000000: data = 6'b000000;
12'b11010101000001: data = 6'b000000;
12'b11010101000010: data = 6'b000000;
12'b11010101000011: data = 6'b000000;
12'b11010101000100: data = 6'b000000;
12'b11010101000101: data = 6'b000000;
12'b11010101000110: data = 6'b000000;
12'b11010101000111: data = 6'b000000;
12'b11010101001000: data = 6'b000000;
12'b11010101001001: data = 6'b000000;
12'b11010101001010: data = 6'b000000;
12'b11010101001011: data = 6'b000000;
12'b11010101001100: data = 6'b000000;
12'b11010101001101: data = 6'b000000;
12'b11010101001110: data = 6'b000000;
12'b11010101001111: data = 6'b000000;
12'b11010101010000: data = 6'b000000;
12'b11010101010001: data = 6'b000000;
12'b11010101010010: data = 6'b000000;
12'b11010101010011: data = 6'b000000;
12'b11010101010100: data = 6'b000000;
12'b11010101010101: data = 6'b000000;
12'b11010101010110: data = 6'b000000;
12'b11010101010111: data = 6'b000000;
12'b11010101011000: data = 6'b000000;
12'b11010101011001: data = 6'b000000;
12'b11010101011010: data = 6'b000000;
12'b11010101011011: data = 6'b000000;
12'b11010101011100: data = 6'b000000;
12'b11010101011101: data = 6'b000000;
12'b11010101011110: data = 6'b000000;
12'b11010101011111: data = 6'b000000;
12'b11010101100000: data = 6'b000000;
12'b11010101100001: data = 6'b000000;
12'b11010101100010: data = 6'b000000;
12'b11010101100011: data = 6'b000000;
12'b11010101100100: data = 6'b000000;
12'b11010101100101: data = 6'b000000;
12'b11010101100110: data = 6'b000000;
12'b11010101100111: data = 6'b000000;
12'b11010101101000: data = 6'b000000;
12'b11010101101001: data = 6'b000000;
12'b11010101101010: data = 6'b000000;
12'b11010101101011: data = 6'b000000;
12'b11010101101100: data = 6'b000000;
12'b11010101101101: data = 6'b000000;
12'b11010101101110: data = 6'b000000;
12'b11010101101111: data = 6'b000000;
12'b11010101110000: data = 6'b000000;
12'b11010101110001: data = 6'b000000;
12'b11010101110010: data = 6'b000000;
12'b11010101110011: data = 6'b000000;
12'b11010101110100: data = 6'b000000;
12'b11010101110101: data = 6'b000000;
12'b11010101110110: data = 6'b000000;
12'b11010101110111: data = 6'b000000;
12'b11010101111000: data = 6'b000000;
12'b11010101111001: data = 6'b000000;
12'b11010101111010: data = 6'b000000;
12'b11010101111011: data = 6'b000000;
12'b11010101111100: data = 6'b000000;
12'b11010101111101: data = 6'b000000;
12'b11010101111110: data = 6'b000000;
12'b11010101111111: data = 6'b000000;
12'b110101010000000: data = 6'b000000;
12'b110101010000001: data = 6'b000000;
12'b110101010000010: data = 6'b000000;
12'b110101010000011: data = 6'b000000;
12'b110101010000100: data = 6'b010101;
12'b110101010000101: data = 6'b010101;
12'b110101010000110: data = 6'b010101;
12'b110101010000111: data = 6'b010101;
12'b110101010001000: data = 6'b010101;
12'b110101010001001: data = 6'b010101;
12'b110101010001010: data = 6'b010101;
12'b110101010001011: data = 6'b010101;
12'b110101010001100: data = 6'b010101;
12'b110101010001101: data = 6'b010101;
12'b110101010001110: data = 6'b101010;
12'b110101010001111: data = 6'b101010;
12'b110101010010000: data = 6'b101010;
12'b110101010010001: data = 6'b101010;
12'b110101010010010: data = 6'b010101;
12'b110101010010011: data = 6'b010101;
12'b110101010010100: data = 6'b010101;
12'b110101010010101: data = 6'b010101;
12'b110101010010110: data = 6'b010101;
12'b110101010010111: data = 6'b010101;
12'b110101010011000: data = 6'b010101;
12'b110101010011001: data = 6'b010101;
12'b110101010011010: data = 6'b010101;
12'b110101010011011: data = 6'b010101;
12'b110101010011100: data = 6'b010101;
12'b110101010011101: data = 6'b010101;
12'b110101010011110: data = 6'b010101;
12'b110101010011111: data = 6'b010101;
12'b110101010100000: data = 6'b010101;
12'b110101010100001: data = 6'b010101;
12'b110101010100010: data = 6'b010101;
12'b110101010100011: data = 6'b010101;
12'b110101010100100: data = 6'b010101;
12'b110101010100101: data = 6'b010101;
12'b110101010100110: data = 6'b010101;
12'b110101010100111: data = 6'b010101;
12'b110101010101000: data = 6'b010101;
12'b110101010101001: data = 6'b010101;
12'b110101010101010: data = 6'b010101;
12'b1101011000000: data = 6'b010101;
12'b1101011000001: data = 6'b010101;
12'b1101011000010: data = 6'b010101;
12'b1101011000011: data = 6'b010101;
12'b1101011000100: data = 6'b010101;
12'b1101011000101: data = 6'b010101;
12'b1101011000110: data = 6'b010101;
12'b1101011000111: data = 6'b010101;
12'b1101011001000: data = 6'b010101;
12'b1101011001001: data = 6'b010101;
12'b1101011001010: data = 6'b010101;
12'b1101011001011: data = 6'b010101;
12'b1101011001100: data = 6'b010101;
12'b1101011001101: data = 6'b010101;
12'b1101011001110: data = 6'b010101;
12'b1101011001111: data = 6'b010101;
12'b1101011010000: data = 6'b010101;
12'b1101011010001: data = 6'b010101;
12'b1101011010010: data = 6'b010101;
12'b1101011010011: data = 6'b010101;
12'b1101011010100: data = 6'b010101;
12'b1101011010101: data = 6'b010101;
12'b1101011010110: data = 6'b010101;
12'b1101011010111: data = 6'b010101;
12'b1101011011000: data = 6'b010101;
12'b1101011011001: data = 6'b101010;
12'b1101011011010: data = 6'b101010;
12'b1101011011011: data = 6'b101010;
12'b1101011011100: data = 6'b101010;
12'b1101011011101: data = 6'b101010;
12'b1101011011110: data = 6'b101010;
12'b1101011011111: data = 6'b101010;
12'b1101011100000: data = 6'b101010;
12'b1101011100001: data = 6'b101010;
12'b1101011100010: data = 6'b010101;
12'b1101011100011: data = 6'b010101;
12'b1101011100100: data = 6'b010101;
12'b1101011100101: data = 6'b010101;
12'b1101011100110: data = 6'b010101;
12'b1101011100111: data = 6'b010101;
12'b1101011101000: data = 6'b010101;
12'b1101011101001: data = 6'b010101;
12'b1101011101010: data = 6'b010101;
12'b1101011101011: data = 6'b010101;
12'b1101011101100: data = 6'b010101;
12'b1101011101101: data = 6'b010101;
12'b1101011101110: data = 6'b010101;
12'b1101011101111: data = 6'b010101;
12'b1101011110000: data = 6'b010101;
12'b1101011110001: data = 6'b010101;
12'b1101011110010: data = 6'b010101;
12'b1101011110011: data = 6'b010101;
12'b1101011110100: data = 6'b010101;
12'b1101011110101: data = 6'b010101;
12'b1101011110110: data = 6'b010101;
12'b1101011110111: data = 6'b010101;
12'b1101011111000: data = 6'b010101;
12'b1101011111001: data = 6'b010101;
12'b1101011111010: data = 6'b010101;
12'b1101011111011: data = 6'b010101;
12'b1101011111100: data = 6'b010101;
12'b1101011111101: data = 6'b010101;
12'b1101011111110: data = 6'b010101;
12'b1101011111111: data = 6'b010101;
12'b11010111000000: data = 6'b010101;
12'b11010111000001: data = 6'b010101;
12'b11010111000010: data = 6'b010101;
12'b11010111000011: data = 6'b010101;
12'b11010111000100: data = 6'b010101;
12'b11010111000101: data = 6'b010101;
12'b11010111000110: data = 6'b010101;
12'b11010111000111: data = 6'b010101;
12'b11010111001000: data = 6'b010101;
12'b11010111001001: data = 6'b010101;
12'b11010111001010: data = 6'b010101;
12'b11010111001011: data = 6'b010101;
12'b11010111001100: data = 6'b010101;
12'b11010111001101: data = 6'b010101;
12'b11010111001110: data = 6'b010101;
12'b11010111001111: data = 6'b010101;
12'b11010111010000: data = 6'b010101;
12'b11010111010001: data = 6'b010101;
12'b11010111010010: data = 6'b010101;
12'b11010111010011: data = 6'b010101;
12'b11010111010100: data = 6'b010101;
12'b11010111010101: data = 6'b010101;
12'b11010111010110: data = 6'b010101;
12'b11010111010111: data = 6'b010101;
12'b11010111011000: data = 6'b010101;
12'b11010111011001: data = 6'b010101;
12'b11010111011010: data = 6'b010101;
12'b11010111011011: data = 6'b010101;
12'b11010111011100: data = 6'b010101;
12'b11010111011101: data = 6'b010101;
12'b11010111011110: data = 6'b010101;
12'b11010111011111: data = 6'b010101;
12'b11010111100000: data = 6'b010101;
12'b11010111100001: data = 6'b010101;
12'b11010111100010: data = 6'b010101;
12'b11010111100011: data = 6'b010101;
12'b11010111100100: data = 6'b010101;
12'b11010111100101: data = 6'b010101;
12'b11010111100110: data = 6'b010101;
12'b11010111100111: data = 6'b010101;
12'b11010111101000: data = 6'b010101;
12'b11010111101001: data = 6'b010101;
12'b11010111101010: data = 6'b010101;
12'b11010111101011: data = 6'b010101;
12'b11010111101100: data = 6'b010101;
12'b11010111101101: data = 6'b010101;
12'b11010111101110: data = 6'b010101;
12'b11010111101111: data = 6'b010101;
12'b11010111110000: data = 6'b010101;
12'b11010111110001: data = 6'b010101;
12'b11010111110010: data = 6'b010101;
12'b11010111110011: data = 6'b010101;
12'b11010111110100: data = 6'b010101;
12'b11010111110101: data = 6'b010101;
12'b11010111110110: data = 6'b010101;
12'b11010111110111: data = 6'b010101;
12'b11010111111000: data = 6'b010101;
12'b11010111111001: data = 6'b010101;
12'b11010111111010: data = 6'b010101;
12'b11010111111011: data = 6'b010101;
12'b11010111111100: data = 6'b010101;
12'b11010111111101: data = 6'b010101;
12'b11010111111110: data = 6'b010101;
12'b11010111111111: data = 6'b010101;
12'b110101110000000: data = 6'b010101;
12'b110101110000001: data = 6'b010101;
12'b110101110000010: data = 6'b010101;
12'b110101110000011: data = 6'b010101;
12'b110101110000100: data = 6'b010101;
12'b110101110000101: data = 6'b010101;
12'b110101110000110: data = 6'b010101;
12'b110101110000111: data = 6'b010101;
12'b110101110001000: data = 6'b010101;
12'b110101110001001: data = 6'b101010;
12'b110101110001010: data = 6'b101010;
12'b110101110001011: data = 6'b101010;
12'b110101110001100: data = 6'b101010;
12'b110101110001101: data = 6'b101010;
12'b110101110001110: data = 6'b101010;
12'b110101110001111: data = 6'b101010;
12'b110101110010000: data = 6'b101010;
12'b110101110010001: data = 6'b101010;
12'b110101110010010: data = 6'b010101;
12'b110101110010011: data = 6'b010101;
12'b110101110010100: data = 6'b010101;
12'b110101110010101: data = 6'b010101;
12'b110101110010110: data = 6'b010101;
12'b110101110010111: data = 6'b010101;
12'b110101110011000: data = 6'b010101;
12'b110101110011001: data = 6'b010101;
12'b110101110011010: data = 6'b010101;
12'b110101110011011: data = 6'b010101;
12'b110101110011100: data = 6'b010101;
12'b110101110011101: data = 6'b010101;
12'b110101110011110: data = 6'b010101;
12'b110101110011111: data = 6'b010101;
12'b110101110100000: data = 6'b010101;
12'b110101110100001: data = 6'b010101;
12'b110101110100010: data = 6'b010101;
12'b110101110100011: data = 6'b010101;
12'b110101110100100: data = 6'b010101;
12'b110101110100101: data = 6'b010101;
12'b110101110100110: data = 6'b010101;
12'b110101110100111: data = 6'b010101;
12'b110101110101000: data = 6'b010101;
12'b110101110101001: data = 6'b010101;
12'b110101110101010: data = 6'b010101;
12'b1101100000000: data = 6'b010101;
12'b1101100000001: data = 6'b010101;
12'b1101100000010: data = 6'b010101;
12'b1101100000011: data = 6'b010101;
12'b1101100000100: data = 6'b010101;
12'b1101100000101: data = 6'b010101;
12'b1101100000110: data = 6'b010101;
12'b1101100000111: data = 6'b010101;
12'b1101100001000: data = 6'b010101;
12'b1101100001001: data = 6'b010101;
12'b1101100001010: data = 6'b010101;
12'b1101100001011: data = 6'b010101;
12'b1101100001100: data = 6'b010101;
12'b1101100001101: data = 6'b010101;
12'b1101100001110: data = 6'b010101;
12'b1101100001111: data = 6'b010101;
12'b1101100010000: data = 6'b010101;
12'b1101100010001: data = 6'b010101;
12'b1101100010010: data = 6'b010101;
12'b1101100010011: data = 6'b010101;
12'b1101100010100: data = 6'b010101;
12'b1101100010101: data = 6'b010101;
12'b1101100010110: data = 6'b010101;
12'b1101100010111: data = 6'b010101;
12'b1101100011000: data = 6'b010101;
12'b1101100011001: data = 6'b101010;
12'b1101100011010: data = 6'b101010;
12'b1101100011011: data = 6'b101010;
12'b1101100011100: data = 6'b101010;
12'b1101100011101: data = 6'b101010;
12'b1101100011110: data = 6'b101010;
12'b1101100011111: data = 6'b101010;
12'b1101100100000: data = 6'b101010;
12'b1101100100001: data = 6'b101010;
12'b1101100100010: data = 6'b010101;
12'b1101100100011: data = 6'b010101;
12'b1101100100100: data = 6'b010101;
12'b1101100100101: data = 6'b010101;
12'b1101100100110: data = 6'b010101;
12'b1101100100111: data = 6'b010101;
12'b1101100101000: data = 6'b010101;
12'b1101100101001: data = 6'b010101;
12'b1101100101010: data = 6'b010101;
12'b1101100101011: data = 6'b010101;
12'b1101100101100: data = 6'b010101;
12'b1101100101101: data = 6'b010101;
12'b1101100101110: data = 6'b010101;
12'b1101100101111: data = 6'b010101;
12'b1101100110000: data = 6'b010101;
12'b1101100110001: data = 6'b010101;
12'b1101100110010: data = 6'b010101;
12'b1101100110011: data = 6'b010101;
12'b1101100110100: data = 6'b010101;
12'b1101100110101: data = 6'b010101;
12'b1101100110110: data = 6'b010101;
12'b1101100110111: data = 6'b010101;
12'b1101100111000: data = 6'b010101;
12'b1101100111001: data = 6'b010101;
12'b1101100111010: data = 6'b010101;
12'b1101100111011: data = 6'b010101;
12'b1101100111100: data = 6'b010101;
12'b1101100111101: data = 6'b010101;
12'b1101100111110: data = 6'b010101;
12'b1101100111111: data = 6'b010101;
12'b11011001000000: data = 6'b010101;
12'b11011001000001: data = 6'b010101;
12'b11011001000010: data = 6'b010101;
12'b11011001000011: data = 6'b010101;
12'b11011001000100: data = 6'b010101;
12'b11011001000101: data = 6'b010101;
12'b11011001000110: data = 6'b010101;
12'b11011001000111: data = 6'b010101;
12'b11011001001000: data = 6'b010101;
12'b11011001001001: data = 6'b010101;
12'b11011001001010: data = 6'b010101;
12'b11011001001011: data = 6'b010101;
12'b11011001001100: data = 6'b010101;
12'b11011001001101: data = 6'b010101;
12'b11011001001110: data = 6'b010101;
12'b11011001001111: data = 6'b010101;
12'b11011001010000: data = 6'b010101;
12'b11011001010001: data = 6'b010101;
12'b11011001010010: data = 6'b010101;
12'b11011001010011: data = 6'b010101;
12'b11011001010100: data = 6'b010101;
12'b11011001010101: data = 6'b010101;
12'b11011001010110: data = 6'b010101;
12'b11011001010111: data = 6'b010101;
12'b11011001011000: data = 6'b010101;
12'b11011001011001: data = 6'b010101;
12'b11011001011010: data = 6'b010101;
12'b11011001011011: data = 6'b010101;
12'b11011001011100: data = 6'b010101;
12'b11011001011101: data = 6'b010101;
12'b11011001011110: data = 6'b010101;
12'b11011001011111: data = 6'b010101;
12'b11011001100000: data = 6'b010101;
12'b11011001100001: data = 6'b010101;
12'b11011001100010: data = 6'b010101;
12'b11011001100011: data = 6'b010101;
12'b11011001100100: data = 6'b010101;
12'b11011001100101: data = 6'b010101;
12'b11011001100110: data = 6'b010101;
12'b11011001100111: data = 6'b010101;
12'b11011001101000: data = 6'b010101;
12'b11011001101001: data = 6'b010101;
12'b11011001101010: data = 6'b010101;
12'b11011001101011: data = 6'b010101;
12'b11011001101100: data = 6'b010101;
12'b11011001101101: data = 6'b010101;
12'b11011001101110: data = 6'b010101;
12'b11011001101111: data = 6'b010101;
12'b11011001110000: data = 6'b010101;
12'b11011001110001: data = 6'b010101;
12'b11011001110010: data = 6'b010101;
12'b11011001110011: data = 6'b010101;
12'b11011001110100: data = 6'b010101;
12'b11011001110101: data = 6'b010101;
12'b11011001110110: data = 6'b010101;
12'b11011001110111: data = 6'b010101;
12'b11011001111000: data = 6'b010101;
12'b11011001111001: data = 6'b010101;
12'b11011001111010: data = 6'b010101;
12'b11011001111011: data = 6'b010101;
12'b11011001111100: data = 6'b010101;
12'b11011001111101: data = 6'b010101;
12'b11011001111110: data = 6'b010101;
12'b11011001111111: data = 6'b010101;
12'b110110010000000: data = 6'b010101;
12'b110110010000001: data = 6'b010101;
12'b110110010000010: data = 6'b010101;
12'b110110010000011: data = 6'b010101;
12'b110110010000100: data = 6'b010101;
12'b110110010000101: data = 6'b010101;
12'b110110010000110: data = 6'b010101;
12'b110110010000111: data = 6'b010101;
12'b110110010001000: data = 6'b010101;
12'b110110010001001: data = 6'b101010;
12'b110110010001010: data = 6'b101010;
12'b110110010001011: data = 6'b101010;
12'b110110010001100: data = 6'b101010;
12'b110110010001101: data = 6'b101010;
12'b110110010001110: data = 6'b101010;
12'b110110010001111: data = 6'b101010;
12'b110110010010000: data = 6'b101010;
12'b110110010010001: data = 6'b101010;
12'b110110010010010: data = 6'b010101;
12'b110110010010011: data = 6'b010101;
12'b110110010010100: data = 6'b010101;
12'b110110010010101: data = 6'b010101;
12'b110110010010110: data = 6'b010101;
12'b110110010010111: data = 6'b010101;
12'b110110010011000: data = 6'b010101;
12'b110110010011001: data = 6'b010101;
12'b110110010011010: data = 6'b010101;
12'b110110010011011: data = 6'b010101;
12'b110110010011100: data = 6'b010101;
12'b110110010011101: data = 6'b010101;
12'b110110010011110: data = 6'b010101;
12'b110110010011111: data = 6'b010101;
12'b110110010100000: data = 6'b010101;
12'b110110010100001: data = 6'b010101;
12'b110110010100010: data = 6'b010101;
12'b110110010100011: data = 6'b010101;
12'b110110010100100: data = 6'b010101;
12'b110110010100101: data = 6'b010101;
12'b110110010100110: data = 6'b010101;
12'b110110010100111: data = 6'b010101;
12'b110110010101000: data = 6'b010101;
12'b110110010101001: data = 6'b010101;
12'b110110010101010: data = 6'b010101;
12'b1101101000000: data = 6'b010101;
12'b1101101000001: data = 6'b010101;
12'b1101101000010: data = 6'b010101;
12'b1101101000011: data = 6'b010101;
12'b1101101000100: data = 6'b010101;
12'b1101101000101: data = 6'b010101;
12'b1101101000110: data = 6'b010101;
12'b1101101000111: data = 6'b010101;
12'b1101101001000: data = 6'b010101;
12'b1101101001001: data = 6'b010101;
12'b1101101001010: data = 6'b010101;
12'b1101101001011: data = 6'b010101;
12'b1101101001100: data = 6'b010101;
12'b1101101001101: data = 6'b010101;
12'b1101101001110: data = 6'b010101;
12'b1101101001111: data = 6'b010101;
12'b1101101010000: data = 6'b010101;
12'b1101101010001: data = 6'b010101;
12'b1101101010010: data = 6'b010101;
12'b1101101010011: data = 6'b010101;
12'b1101101010100: data = 6'b010101;
12'b1101101010101: data = 6'b010101;
12'b1101101010110: data = 6'b010101;
12'b1101101010111: data = 6'b010101;
12'b1101101011000: data = 6'b010101;
12'b1101101011001: data = 6'b101010;
12'b1101101011010: data = 6'b101010;
12'b1101101011011: data = 6'b101010;
12'b1101101011100: data = 6'b101010;
12'b1101101011101: data = 6'b101010;
12'b1101101011110: data = 6'b101010;
12'b1101101011111: data = 6'b101010;
12'b1101101100000: data = 6'b101010;
12'b1101101100001: data = 6'b101010;
12'b1101101100010: data = 6'b101010;
12'b1101101100011: data = 6'b101010;
12'b1101101100100: data = 6'b101001;
12'b1101101100101: data = 6'b010101;
12'b1101101100110: data = 6'b010101;
12'b1101101100111: data = 6'b010101;
12'b1101101101000: data = 6'b010101;
12'b1101101101001: data = 6'b010101;
12'b1101101101010: data = 6'b010101;
12'b1101101101011: data = 6'b010101;
12'b1101101101100: data = 6'b010101;
12'b1101101101101: data = 6'b010101;
12'b1101101101110: data = 6'b010101;
12'b1101101101111: data = 6'b010101;
12'b1101101110000: data = 6'b010101;
12'b1101101110001: data = 6'b010101;
12'b1101101110010: data = 6'b010101;
12'b1101101110011: data = 6'b010101;
12'b1101101110100: data = 6'b010101;
12'b1101101110101: data = 6'b010101;
12'b1101101110110: data = 6'b010101;
12'b1101101110111: data = 6'b010101;
12'b1101101111000: data = 6'b010101;
12'b1101101111001: data = 6'b010101;
12'b1101101111010: data = 6'b010101;
12'b1101101111011: data = 6'b010101;
12'b1101101111100: data = 6'b010101;
12'b1101101111101: data = 6'b010101;
12'b1101101111110: data = 6'b010101;
12'b1101101111111: data = 6'b010101;
12'b11011011000000: data = 6'b010101;
12'b11011011000001: data = 6'b010101;
12'b11011011000010: data = 6'b010101;
12'b11011011000011: data = 6'b010101;
12'b11011011000100: data = 6'b010101;
12'b11011011000101: data = 6'b010101;
12'b11011011000110: data = 6'b010101;
12'b11011011000111: data = 6'b010101;
12'b11011011001000: data = 6'b010101;
12'b11011011001001: data = 6'b010101;
12'b11011011001010: data = 6'b010101;
12'b11011011001011: data = 6'b010101;
12'b11011011001100: data = 6'b010101;
12'b11011011001101: data = 6'b010101;
12'b11011011001110: data = 6'b010101;
12'b11011011001111: data = 6'b010101;
12'b11011011010000: data = 6'b010101;
12'b11011011010001: data = 6'b010101;
12'b11011011010010: data = 6'b010101;
12'b11011011010011: data = 6'b010101;
12'b11011011010100: data = 6'b010101;
12'b11011011010101: data = 6'b010101;
12'b11011011010110: data = 6'b010101;
12'b11011011010111: data = 6'b010101;
12'b11011011011000: data = 6'b010101;
12'b11011011011001: data = 6'b010101;
12'b11011011011010: data = 6'b010101;
12'b11011011011011: data = 6'b010101;
12'b11011011011100: data = 6'b010101;
12'b11011011011101: data = 6'b010101;
12'b11011011011110: data = 6'b010101;
12'b11011011011111: data = 6'b010101;
12'b11011011100000: data = 6'b010101;
12'b11011011100001: data = 6'b010101;
12'b11011011100010: data = 6'b010101;
12'b11011011100011: data = 6'b010101;
12'b11011011100100: data = 6'b010101;
12'b11011011100101: data = 6'b010101;
12'b11011011100110: data = 6'b010101;
12'b11011011100111: data = 6'b010101;
12'b11011011101000: data = 6'b010101;
12'b11011011101001: data = 6'b010101;
12'b11011011101010: data = 6'b010101;
12'b11011011101011: data = 6'b010101;
12'b11011011101100: data = 6'b010101;
12'b11011011101101: data = 6'b010101;
12'b11011011101110: data = 6'b010101;
12'b11011011101111: data = 6'b010101;
12'b11011011110000: data = 6'b010101;
12'b11011011110001: data = 6'b010101;
12'b11011011110010: data = 6'b010101;
12'b11011011110011: data = 6'b010101;
12'b11011011110100: data = 6'b010101;
12'b11011011110101: data = 6'b010101;
12'b11011011110110: data = 6'b010101;
12'b11011011110111: data = 6'b010101;
12'b11011011111000: data = 6'b010101;
12'b11011011111001: data = 6'b010101;
12'b11011011111010: data = 6'b010101;
12'b11011011111011: data = 6'b010101;
12'b11011011111100: data = 6'b010101;
12'b11011011111101: data = 6'b010101;
12'b11011011111110: data = 6'b010101;
12'b11011011111111: data = 6'b010101;
12'b110110110000000: data = 6'b010101;
12'b110110110000001: data = 6'b010101;
12'b110110110000010: data = 6'b010101;
12'b110110110000011: data = 6'b010101;
12'b110110110000100: data = 6'b010101;
12'b110110110000101: data = 6'b010101;
12'b110110110000110: data = 6'b010101;
12'b110110110000111: data = 6'b010101;
12'b110110110001000: data = 6'b101010;
12'b110110110001001: data = 6'b101010;
12'b110110110001010: data = 6'b101010;
12'b110110110001011: data = 6'b101010;
12'b110110110001100: data = 6'b101010;
12'b110110110001101: data = 6'b101010;
12'b110110110001110: data = 6'b101010;
12'b110110110001111: data = 6'b101010;
12'b110110110010000: data = 6'b101010;
12'b110110110010001: data = 6'b101010;
12'b110110110010010: data = 6'b010101;
12'b110110110010011: data = 6'b010101;
12'b110110110010100: data = 6'b010101;
12'b110110110010101: data = 6'b010101;
12'b110110110010110: data = 6'b010101;
12'b110110110010111: data = 6'b010101;
12'b110110110011000: data = 6'b010101;
12'b110110110011001: data = 6'b010101;
12'b110110110011010: data = 6'b010101;
12'b110110110011011: data = 6'b010101;
12'b110110110011100: data = 6'b010101;
12'b110110110011101: data = 6'b010101;
12'b110110110011110: data = 6'b010101;
12'b110110110011111: data = 6'b010101;
12'b110110110100000: data = 6'b010101;
12'b110110110100001: data = 6'b010101;
12'b110110110100010: data = 6'b010101;
12'b110110110100011: data = 6'b010101;
12'b110110110100100: data = 6'b010101;
12'b110110110100101: data = 6'b010101;
12'b110110110100110: data = 6'b010101;
12'b110110110100111: data = 6'b010101;
12'b110110110101000: data = 6'b010101;
12'b110110110101001: data = 6'b010101;
12'b110110110101010: data = 6'b010101;
12'b1101110000000: data = 6'b010101;
12'b1101110000001: data = 6'b010101;
12'b1101110000010: data = 6'b010101;
12'b1101110000011: data = 6'b010101;
12'b1101110000100: data = 6'b010101;
12'b1101110000101: data = 6'b010101;
12'b1101110000110: data = 6'b010101;
12'b1101110000111: data = 6'b010101;
12'b1101110001000: data = 6'b010101;
12'b1101110001001: data = 6'b010101;
12'b1101110001010: data = 6'b010101;
12'b1101110001011: data = 6'b010101;
12'b1101110001100: data = 6'b010101;
12'b1101110001101: data = 6'b010101;
12'b1101110001110: data = 6'b010101;
12'b1101110001111: data = 6'b010101;
12'b1101110010000: data = 6'b010101;
12'b1101110010001: data = 6'b010101;
12'b1101110010010: data = 6'b010101;
12'b1101110010011: data = 6'b010101;
12'b1101110010100: data = 6'b010101;
12'b1101110010101: data = 6'b010101;
12'b1101110010110: data = 6'b010101;
12'b1101110010111: data = 6'b010101;
12'b1101110011000: data = 6'b010101;
12'b1101110011001: data = 6'b101010;
12'b1101110011010: data = 6'b101010;
12'b1101110011011: data = 6'b101010;
12'b1101110011100: data = 6'b101010;
12'b1101110011101: data = 6'b101010;
12'b1101110011110: data = 6'b101010;
12'b1101110011111: data = 6'b101010;
12'b1101110100000: data = 6'b101010;
12'b1101110100001: data = 6'b101010;
12'b1101110100010: data = 6'b101010;
12'b1101110100011: data = 6'b101010;
12'b1101110100100: data = 6'b101010;
12'b1101110100101: data = 6'b010101;
12'b1101110100110: data = 6'b010101;
12'b1101110100111: data = 6'b010101;
12'b1101110101000: data = 6'b010101;
12'b1101110101001: data = 6'b010101;
12'b1101110101010: data = 6'b010101;
12'b1101110101011: data = 6'b010101;
12'b1101110101100: data = 6'b010101;
12'b1101110101101: data = 6'b010101;
12'b1101110101110: data = 6'b010101;
12'b1101110101111: data = 6'b010101;
12'b1101110110000: data = 6'b010101;
12'b1101110110001: data = 6'b010101;
12'b1101110110010: data = 6'b010101;
12'b1101110110011: data = 6'b010101;
12'b1101110110100: data = 6'b010101;
12'b1101110110101: data = 6'b010101;
12'b1101110110110: data = 6'b010101;
12'b1101110110111: data = 6'b010101;
12'b1101110111000: data = 6'b010101;
12'b1101110111001: data = 6'b010101;
12'b1101110111010: data = 6'b010101;
12'b1101110111011: data = 6'b010101;
12'b1101110111100: data = 6'b010101;
12'b1101110111101: data = 6'b010101;
12'b1101110111110: data = 6'b010101;
12'b1101110111111: data = 6'b010101;
12'b11011101000000: data = 6'b010101;
12'b11011101000001: data = 6'b010101;
12'b11011101000010: data = 6'b010101;
12'b11011101000011: data = 6'b010101;
12'b11011101000100: data = 6'b010101;
12'b11011101000101: data = 6'b010101;
12'b11011101000110: data = 6'b010101;
12'b11011101000111: data = 6'b010101;
12'b11011101001000: data = 6'b010101;
12'b11011101001001: data = 6'b010101;
12'b11011101001010: data = 6'b010101;
12'b11011101001011: data = 6'b010101;
12'b11011101001100: data = 6'b010101;
12'b11011101001101: data = 6'b010101;
12'b11011101001110: data = 6'b010101;
12'b11011101001111: data = 6'b010101;
12'b11011101010000: data = 6'b010101;
12'b11011101010001: data = 6'b010101;
12'b11011101010010: data = 6'b010101;
12'b11011101010011: data = 6'b010101;
12'b11011101010100: data = 6'b010101;
12'b11011101010101: data = 6'b010101;
12'b11011101010110: data = 6'b010101;
12'b11011101010111: data = 6'b010101;
12'b11011101011000: data = 6'b010101;
12'b11011101011001: data = 6'b010101;
12'b11011101011010: data = 6'b010101;
12'b11011101011011: data = 6'b010101;
12'b11011101011100: data = 6'b010101;
12'b11011101011101: data = 6'b010101;
12'b11011101011110: data = 6'b010101;
12'b11011101011111: data = 6'b010101;
12'b11011101100000: data = 6'b010101;
12'b11011101100001: data = 6'b010101;
12'b11011101100010: data = 6'b010101;
12'b11011101100011: data = 6'b010101;
12'b11011101100100: data = 6'b010101;
12'b11011101100101: data = 6'b010101;
12'b11011101100110: data = 6'b010101;
12'b11011101100111: data = 6'b010101;
12'b11011101101000: data = 6'b010101;
12'b11011101101001: data = 6'b010101;
12'b11011101101010: data = 6'b010101;
12'b11011101101011: data = 6'b010101;
12'b11011101101100: data = 6'b010101;
12'b11011101101101: data = 6'b010101;
12'b11011101101110: data = 6'b010101;
12'b11011101101111: data = 6'b010101;
12'b11011101110000: data = 6'b010101;
12'b11011101110001: data = 6'b010101;
12'b11011101110010: data = 6'b010101;
12'b11011101110011: data = 6'b010101;
12'b11011101110100: data = 6'b010101;
12'b11011101110101: data = 6'b010101;
12'b11011101110110: data = 6'b010101;
12'b11011101110111: data = 6'b010101;
12'b11011101111000: data = 6'b010101;
12'b11011101111001: data = 6'b010101;
12'b11011101111010: data = 6'b010101;
12'b11011101111011: data = 6'b010101;
12'b11011101111100: data = 6'b010101;
12'b11011101111101: data = 6'b010101;
12'b11011101111110: data = 6'b010101;
12'b11011101111111: data = 6'b010101;
12'b110111010000000: data = 6'b010101;
12'b110111010000001: data = 6'b010101;
12'b110111010000010: data = 6'b010101;
12'b110111010000011: data = 6'b010101;
12'b110111010000100: data = 6'b010101;
12'b110111010000101: data = 6'b010101;
12'b110111010000110: data = 6'b101001;
12'b110111010000111: data = 6'b101010;
12'b110111010001000: data = 6'b101010;
12'b110111010001001: data = 6'b101010;
12'b110111010001010: data = 6'b101010;
12'b110111010001011: data = 6'b101010;
12'b110111010001100: data = 6'b101010;
12'b110111010001101: data = 6'b101010;
12'b110111010001110: data = 6'b101010;
12'b110111010001111: data = 6'b101010;
12'b110111010010000: data = 6'b101010;
12'b110111010010001: data = 6'b101010;
12'b110111010010010: data = 6'b010101;
12'b110111010010011: data = 6'b010101;
12'b110111010010100: data = 6'b010101;
12'b110111010010101: data = 6'b010101;
12'b110111010010110: data = 6'b010101;
12'b110111010010111: data = 6'b010101;
12'b110111010011000: data = 6'b010101;
12'b110111010011001: data = 6'b010101;
12'b110111010011010: data = 6'b010101;
12'b110111010011011: data = 6'b010101;
12'b110111010011100: data = 6'b010101;
12'b110111010011101: data = 6'b010101;
12'b110111010011110: data = 6'b010101;
12'b110111010011111: data = 6'b010101;
12'b110111010100000: data = 6'b010101;
12'b110111010100001: data = 6'b010101;
12'b110111010100010: data = 6'b010101;
12'b110111010100011: data = 6'b010101;
12'b110111010100100: data = 6'b010101;
12'b110111010100101: data = 6'b010101;
12'b110111010100110: data = 6'b010101;
12'b110111010100111: data = 6'b010101;
12'b110111010101000: data = 6'b010101;
12'b110111010101001: data = 6'b010101;
12'b110111010101010: data = 6'b010101;
12'b1101111000000: data = 6'b010101;
12'b1101111000001: data = 6'b010101;
12'b1101111000010: data = 6'b010101;
12'b1101111000011: data = 6'b010101;
12'b1101111000100: data = 6'b010101;
12'b1101111000101: data = 6'b010101;
12'b1101111000110: data = 6'b010101;
12'b1101111000111: data = 6'b010101;
12'b1101111001000: data = 6'b010101;
12'b1101111001001: data = 6'b010101;
12'b1101111001010: data = 6'b010101;
12'b1101111001011: data = 6'b010101;
12'b1101111001100: data = 6'b010101;
12'b1101111001101: data = 6'b010101;
12'b1101111001110: data = 6'b010101;
12'b1101111001111: data = 6'b010101;
12'b1101111010000: data = 6'b010101;
12'b1101111010001: data = 6'b010101;
12'b1101111010010: data = 6'b010101;
12'b1101111010011: data = 6'b010101;
12'b1101111010100: data = 6'b010101;
12'b1101111010101: data = 6'b010101;
12'b1101111010110: data = 6'b010101;
12'b1101111010111: data = 6'b010101;
12'b1101111011000: data = 6'b010101;
12'b1101111011001: data = 6'b101010;
12'b1101111011010: data = 6'b101010;
12'b1101111011011: data = 6'b101010;
12'b1101111011100: data = 6'b101010;
12'b1101111011101: data = 6'b101010;
12'b1101111011110: data = 6'b101010;
12'b1101111011111: data = 6'b101010;
12'b1101111100000: data = 6'b101010;
12'b1101111100001: data = 6'b101010;
12'b1101111100010: data = 6'b101010;
12'b1101111100011: data = 6'b101010;
12'b1101111100100: data = 6'b101001;
12'b1101111100101: data = 6'b010101;
12'b1101111100110: data = 6'b010101;
12'b1101111100111: data = 6'b010101;
12'b1101111101000: data = 6'b010101;
12'b1101111101001: data = 6'b010101;
12'b1101111101010: data = 6'b010101;
12'b1101111101011: data = 6'b010101;
12'b1101111101100: data = 6'b010101;
12'b1101111101101: data = 6'b010101;
12'b1101111101110: data = 6'b010101;
12'b1101111101111: data = 6'b010101;
12'b1101111110000: data = 6'b010101;
12'b1101111110001: data = 6'b010101;
12'b1101111110010: data = 6'b010101;
12'b1101111110011: data = 6'b010101;
12'b1101111110100: data = 6'b010101;
12'b1101111110101: data = 6'b010101;
12'b1101111110110: data = 6'b010101;
12'b1101111110111: data = 6'b010101;
12'b1101111111000: data = 6'b010101;
12'b1101111111001: data = 6'b010101;
12'b1101111111010: data = 6'b010101;
12'b1101111111011: data = 6'b010101;
12'b1101111111100: data = 6'b010101;
12'b1101111111101: data = 6'b010101;
12'b1101111111110: data = 6'b010101;
12'b1101111111111: data = 6'b010101;
12'b11011111000000: data = 6'b010101;
12'b11011111000001: data = 6'b010101;
12'b11011111000010: data = 6'b010101;
12'b11011111000011: data = 6'b010101;
12'b11011111000100: data = 6'b010101;
12'b11011111000101: data = 6'b010101;
12'b11011111000110: data = 6'b010101;
12'b11011111000111: data = 6'b010101;
12'b11011111001000: data = 6'b010101;
12'b11011111001001: data = 6'b010101;
12'b11011111001010: data = 6'b010101;
12'b11011111001011: data = 6'b010101;
12'b11011111001100: data = 6'b010101;
12'b11011111001101: data = 6'b010101;
12'b11011111001110: data = 6'b010101;
12'b11011111001111: data = 6'b010101;
12'b11011111010000: data = 6'b010101;
12'b11011111010001: data = 6'b010101;
12'b11011111010010: data = 6'b010101;
12'b11011111010011: data = 6'b010101;
12'b11011111010100: data = 6'b010101;
12'b11011111010101: data = 6'b010101;
12'b11011111010110: data = 6'b010101;
12'b11011111010111: data = 6'b010101;
12'b11011111011000: data = 6'b010101;
12'b11011111011001: data = 6'b010101;
12'b11011111011010: data = 6'b010101;
12'b11011111011011: data = 6'b010101;
12'b11011111011100: data = 6'b010101;
12'b11011111011101: data = 6'b010101;
12'b11011111011110: data = 6'b010101;
12'b11011111011111: data = 6'b010101;
12'b11011111100000: data = 6'b010101;
12'b11011111100001: data = 6'b010101;
12'b11011111100010: data = 6'b010101;
12'b11011111100011: data = 6'b010101;
12'b11011111100100: data = 6'b010101;
12'b11011111100101: data = 6'b010101;
12'b11011111100110: data = 6'b010101;
12'b11011111100111: data = 6'b010101;
12'b11011111101000: data = 6'b010101;
12'b11011111101001: data = 6'b010101;
12'b11011111101010: data = 6'b010101;
12'b11011111101011: data = 6'b010101;
12'b11011111101100: data = 6'b010101;
12'b11011111101101: data = 6'b010101;
12'b11011111101110: data = 6'b010101;
12'b11011111101111: data = 6'b010101;
12'b11011111110000: data = 6'b010101;
12'b11011111110001: data = 6'b010101;
12'b11011111110010: data = 6'b010101;
12'b11011111110011: data = 6'b010101;
12'b11011111110100: data = 6'b010101;
12'b11011111110101: data = 6'b010101;
12'b11011111110110: data = 6'b010101;
12'b11011111110111: data = 6'b010101;
12'b11011111111000: data = 6'b010101;
12'b11011111111001: data = 6'b010101;
12'b11011111111010: data = 6'b010101;
12'b11011111111011: data = 6'b010101;
12'b11011111111100: data = 6'b010101;
12'b11011111111101: data = 6'b010101;
12'b11011111111110: data = 6'b010101;
12'b11011111111111: data = 6'b010101;
12'b110111110000000: data = 6'b010101;
12'b110111110000001: data = 6'b010101;
12'b110111110000010: data = 6'b010101;
12'b110111110000011: data = 6'b010101;
12'b110111110000100: data = 6'b010101;
12'b110111110000101: data = 6'b010101;
12'b110111110000110: data = 6'b010101;
12'b110111110000111: data = 6'b101001;
12'b110111110001000: data = 6'b101010;
12'b110111110001001: data = 6'b101010;
12'b110111110001010: data = 6'b101010;
12'b110111110001011: data = 6'b101010;
12'b110111110001100: data = 6'b101010;
12'b110111110001101: data = 6'b101010;
12'b110111110001110: data = 6'b101010;
12'b110111110001111: data = 6'b101010;
12'b110111110010000: data = 6'b101010;
12'b110111110010001: data = 6'b101010;
12'b110111110010010: data = 6'b010101;
12'b110111110010011: data = 6'b010101;
12'b110111110010100: data = 6'b010101;
12'b110111110010101: data = 6'b010101;
12'b110111110010110: data = 6'b010101;
12'b110111110010111: data = 6'b010101;
12'b110111110011000: data = 6'b010101;
12'b110111110011001: data = 6'b010101;
12'b110111110011010: data = 6'b010101;
12'b110111110011011: data = 6'b010101;
12'b110111110011100: data = 6'b010101;
12'b110111110011101: data = 6'b010101;
12'b110111110011110: data = 6'b010101;
12'b110111110011111: data = 6'b010101;
12'b110111110100000: data = 6'b010101;
12'b110111110100001: data = 6'b010101;
12'b110111110100010: data = 6'b010101;
12'b110111110100011: data = 6'b010101;
12'b110111110100100: data = 6'b010101;
12'b110111110100101: data = 6'b010101;
12'b110111110100110: data = 6'b010101;
12'b110111110100111: data = 6'b010101;
12'b110111110101000: data = 6'b010101;
12'b110111110101001: data = 6'b010101;
12'b110111110101010: data = 6'b010101;
12'b1110000000000: data = 6'b010101;
12'b1110000000001: data = 6'b010101;
12'b1110000000010: data = 6'b010101;
12'b1110000000011: data = 6'b010101;
12'b1110000000100: data = 6'b010101;
12'b1110000000101: data = 6'b010101;
12'b1110000000110: data = 6'b010101;
12'b1110000000111: data = 6'b010101;
12'b1110000001000: data = 6'b010101;
12'b1110000001001: data = 6'b010101;
12'b1110000001010: data = 6'b010101;
12'b1110000001011: data = 6'b010101;
12'b1110000001100: data = 6'b010101;
12'b1110000001101: data = 6'b010101;
12'b1110000001110: data = 6'b010101;
12'b1110000001111: data = 6'b010101;
12'b1110000010000: data = 6'b010101;
12'b1110000010001: data = 6'b010101;
12'b1110000010010: data = 6'b010101;
12'b1110000010011: data = 6'b010101;
12'b1110000010100: data = 6'b010101;
12'b1110000010101: data = 6'b010101;
12'b1110000010110: data = 6'b010101;
12'b1110000010111: data = 6'b010101;
12'b1110000011000: data = 6'b010101;
12'b1110000011001: data = 6'b101010;
12'b1110000011010: data = 6'b101010;
12'b1110000011011: data = 6'b101010;
12'b1110000011100: data = 6'b101001;
12'b1110000011101: data = 6'b010101;
12'b1110000011110: data = 6'b000000;
12'b1110000011111: data = 6'b000000;
12'b1110000100000: data = 6'b000000;
12'b1110000100001: data = 6'b000000;
12'b1110000100010: data = 6'b000000;
12'b1110000100011: data = 6'b000000;
12'b1110000100100: data = 6'b000000;
12'b1110000100101: data = 6'b000000;
12'b1110000100110: data = 6'b000000;
12'b1110000100111: data = 6'b000000;
12'b1110000101000: data = 6'b000000;
12'b1110000101001: data = 6'b000000;
12'b1110000101010: data = 6'b000000;
12'b1110000101011: data = 6'b000000;
12'b1110000101100: data = 6'b000000;
12'b1110000101101: data = 6'b000000;
12'b1110000101110: data = 6'b000000;
12'b1110000101111: data = 6'b010101;
12'b1110000110000: data = 6'b010101;
12'b1110000110001: data = 6'b010101;
12'b1110000110010: data = 6'b010101;
12'b1110000110011: data = 6'b010101;
12'b1110000110100: data = 6'b010101;
12'b1110000110101: data = 6'b010101;
12'b1110000110110: data = 6'b010101;
12'b1110000110111: data = 6'b010101;
12'b1110000111000: data = 6'b010101;
12'b1110000111001: data = 6'b010101;
12'b1110000111010: data = 6'b010101;
12'b1110000111011: data = 6'b010101;
12'b1110000111100: data = 6'b010101;
12'b1110000111101: data = 6'b010101;
12'b1110000111110: data = 6'b010101;
12'b1110000111111: data = 6'b010101;
12'b11100001000000: data = 6'b010101;
12'b11100001000001: data = 6'b010101;
12'b11100001000010: data = 6'b010101;
12'b11100001000011: data = 6'b010101;
12'b11100001000100: data = 6'b010101;
12'b11100001000101: data = 6'b010101;
12'b11100001000110: data = 6'b010101;
12'b11100001000111: data = 6'b010101;
12'b11100001001000: data = 6'b010101;
12'b11100001001001: data = 6'b010101;
12'b11100001001010: data = 6'b010101;
12'b11100001001011: data = 6'b010101;
12'b11100001001100: data = 6'b010101;
12'b11100001001101: data = 6'b010101;
12'b11100001001110: data = 6'b010101;
12'b11100001001111: data = 6'b010101;
12'b11100001010000: data = 6'b010101;
12'b11100001010001: data = 6'b010101;
12'b11100001010010: data = 6'b010101;
12'b11100001010011: data = 6'b010101;
12'b11100001010100: data = 6'b010101;
12'b11100001010101: data = 6'b010101;
12'b11100001010110: data = 6'b010101;
12'b11100001010111: data = 6'b010101;
12'b11100001011000: data = 6'b010101;
12'b11100001011001: data = 6'b010101;
12'b11100001011010: data = 6'b010101;
12'b11100001011011: data = 6'b010101;
12'b11100001011100: data = 6'b010101;
12'b11100001011101: data = 6'b010101;
12'b11100001011110: data = 6'b010101;
12'b11100001011111: data = 6'b010101;
12'b11100001100000: data = 6'b010101;
12'b11100001100001: data = 6'b010101;
12'b11100001100010: data = 6'b010101;
12'b11100001100011: data = 6'b010101;
12'b11100001100100: data = 6'b010101;
12'b11100001100101: data = 6'b010101;
12'b11100001100110: data = 6'b010101;
12'b11100001100111: data = 6'b010101;
12'b11100001101000: data = 6'b010101;
12'b11100001101001: data = 6'b010101;
12'b11100001101010: data = 6'b010101;
12'b11100001101011: data = 6'b010101;
12'b11100001101100: data = 6'b010101;
12'b11100001101101: data = 6'b010101;
12'b11100001101110: data = 6'b010101;
12'b11100001101111: data = 6'b010101;
12'b11100001110000: data = 6'b010101;
12'b11100001110001: data = 6'b010101;
12'b11100001110010: data = 6'b010101;
12'b11100001110011: data = 6'b010101;
12'b11100001110100: data = 6'b010101;
12'b11100001110101: data = 6'b010101;
12'b11100001110110: data = 6'b010101;
12'b11100001110111: data = 6'b010101;
12'b11100001111000: data = 6'b010101;
12'b11100001111001: data = 6'b010101;
12'b11100001111010: data = 6'b010101;
12'b11100001111011: data = 6'b010101;
12'b11100001111100: data = 6'b010101;
12'b11100001111101: data = 6'b010101;
12'b11100001111110: data = 6'b010101;
12'b11100001111111: data = 6'b010101;
12'b111000010000000: data = 6'b000000;
12'b111000010000001: data = 6'b000000;
12'b111000010000010: data = 6'b000000;
12'b111000010000011: data = 6'b000000;
12'b111000010000100: data = 6'b000000;
12'b111000010000101: data = 6'b000000;
12'b111000010000110: data = 6'b000000;
12'b111000010000111: data = 6'b000000;
12'b111000010001000: data = 6'b000000;
12'b111000010001001: data = 6'b000000;
12'b111000010001010: data = 6'b000000;
12'b111000010001011: data = 6'b010101;
12'b111000010001100: data = 6'b010101;
12'b111000010001101: data = 6'b010101;
12'b111000010001110: data = 6'b101010;
12'b111000010001111: data = 6'b101010;
12'b111000010010000: data = 6'b101010;
12'b111000010010001: data = 6'b101010;
12'b111000010010010: data = 6'b010101;
12'b111000010010011: data = 6'b010101;
12'b111000010010100: data = 6'b010101;
12'b111000010010101: data = 6'b010101;
12'b111000010010110: data = 6'b010101;
12'b111000010010111: data = 6'b010101;
12'b111000010011000: data = 6'b010101;
12'b111000010011001: data = 6'b010101;
12'b111000010011010: data = 6'b010101;
12'b111000010011011: data = 6'b010101;
12'b111000010011100: data = 6'b010101;
12'b111000010011101: data = 6'b010101;
12'b111000010011110: data = 6'b010101;
12'b111000010011111: data = 6'b010101;
12'b111000010100000: data = 6'b010101;
12'b111000010100001: data = 6'b010101;
12'b111000010100010: data = 6'b010101;
12'b111000010100011: data = 6'b010101;
12'b111000010100100: data = 6'b010101;
12'b111000010100101: data = 6'b010101;
12'b111000010100110: data = 6'b010101;
12'b111000010100111: data = 6'b010101;
12'b111000010101000: data = 6'b010101;
12'b111000010101001: data = 6'b010101;
12'b111000010101010: data = 6'b010101;
12'b1110001000000: data = 6'b010101;
12'b1110001000001: data = 6'b010101;
12'b1110001000010: data = 6'b010101;
12'b1110001000011: data = 6'b010101;
12'b1110001000100: data = 6'b010101;
12'b1110001000101: data = 6'b010101;
12'b1110001000110: data = 6'b010101;
12'b1110001000111: data = 6'b010101;
12'b1110001001000: data = 6'b010101;
12'b1110001001001: data = 6'b010101;
12'b1110001001010: data = 6'b010101;
12'b1110001001011: data = 6'b010101;
12'b1110001001100: data = 6'b010101;
12'b1110001001101: data = 6'b010101;
12'b1110001001110: data = 6'b010101;
12'b1110001001111: data = 6'b010101;
12'b1110001010000: data = 6'b010101;
12'b1110001010001: data = 6'b010101;
12'b1110001010010: data = 6'b010101;
12'b1110001010011: data = 6'b010101;
12'b1110001010100: data = 6'b010101;
12'b1110001010101: data = 6'b010101;
12'b1110001010110: data = 6'b010101;
12'b1110001010111: data = 6'b010101;
12'b1110001011000: data = 6'b010101;
12'b1110001011001: data = 6'b101010;
12'b1110001011010: data = 6'b101010;
12'b1110001011011: data = 6'b101010;
12'b1110001011100: data = 6'b010101;
12'b1110001011101: data = 6'b000000;
12'b1110001011110: data = 6'b000000;
12'b1110001011111: data = 6'b000000;
12'b1110001100000: data = 6'b000000;
12'b1110001100001: data = 6'b000000;
12'b1110001100010: data = 6'b000000;
12'b1110001100011: data = 6'b000000;
12'b1110001100100: data = 6'b000000;
12'b1110001100101: data = 6'b000000;
12'b1110001100110: data = 6'b000000;
12'b1110001100111: data = 6'b000000;
12'b1110001101000: data = 6'b000000;
12'b1110001101001: data = 6'b000000;
12'b1110001101010: data = 6'b000000;
12'b1110001101011: data = 6'b000000;
12'b1110001101100: data = 6'b000000;
12'b1110001101101: data = 6'b000000;
12'b1110001101110: data = 6'b000000;
12'b1110001101111: data = 6'b000000;
12'b1110001110000: data = 6'b000000;
12'b1110001110001: data = 6'b000000;
12'b1110001110010: data = 6'b000000;
12'b1110001110011: data = 6'b000000;
12'b1110001110100: data = 6'b000000;
12'b1110001110101: data = 6'b010101;
12'b1110001110110: data = 6'b000000;
12'b1110001110111: data = 6'b010101;
12'b1110001111000: data = 6'b010101;
12'b1110001111001: data = 6'b010101;
12'b1110001111010: data = 6'b010101;
12'b1110001111011: data = 6'b010101;
12'b1110001111100: data = 6'b010101;
12'b1110001111101: data = 6'b010101;
12'b1110001111110: data = 6'b010101;
12'b1110001111111: data = 6'b010101;
12'b11100011000000: data = 6'b010101;
12'b11100011000001: data = 6'b010101;
12'b11100011000010: data = 6'b010101;
12'b11100011000011: data = 6'b010101;
12'b11100011000100: data = 6'b010101;
12'b11100011000101: data = 6'b010101;
12'b11100011000110: data = 6'b010101;
12'b11100011000111: data = 6'b010101;
12'b11100011001000: data = 6'b010101;
12'b11100011001001: data = 6'b010101;
12'b11100011001010: data = 6'b010101;
12'b11100011001011: data = 6'b010101;
12'b11100011001100: data = 6'b010101;
12'b11100011001101: data = 6'b010101;
12'b11100011001110: data = 6'b010101;
12'b11100011001111: data = 6'b010101;
12'b11100011010000: data = 6'b010101;
12'b11100011010001: data = 6'b010101;
12'b11100011010010: data = 6'b010101;
12'b11100011010011: data = 6'b010101;
12'b11100011010100: data = 6'b010101;
12'b11100011010101: data = 6'b010101;
12'b11100011010110: data = 6'b010101;
12'b11100011010111: data = 6'b010101;
12'b11100011011000: data = 6'b010101;
12'b11100011011001: data = 6'b010101;
12'b11100011011010: data = 6'b010101;
12'b11100011011011: data = 6'b010101;
12'b11100011011100: data = 6'b010101;
12'b11100011011101: data = 6'b010101;
12'b11100011011110: data = 6'b010101;
12'b11100011011111: data = 6'b010101;
12'b11100011100000: data = 6'b010101;
12'b11100011100001: data = 6'b010101;
12'b11100011100010: data = 6'b010101;
12'b11100011100011: data = 6'b010101;
12'b11100011100100: data = 6'b010101;
12'b11100011100101: data = 6'b010101;
12'b11100011100110: data = 6'b010101;
12'b11100011100111: data = 6'b010101;
12'b11100011101000: data = 6'b010101;
12'b11100011101001: data = 6'b010101;
12'b11100011101010: data = 6'b010101;
12'b11100011101011: data = 6'b010101;
12'b11100011101100: data = 6'b010101;
12'b11100011101101: data = 6'b010101;
12'b11100011101110: data = 6'b010101;
12'b11100011101111: data = 6'b010101;
12'b11100011110000: data = 6'b010101;
12'b11100011110001: data = 6'b010101;
12'b11100011110010: data = 6'b010101;
12'b11100011110011: data = 6'b010101;
12'b11100011110100: data = 6'b010101;
12'b11100011110101: data = 6'b010101;
12'b11100011110110: data = 6'b010101;
12'b11100011110111: data = 6'b000000;
12'b11100011111000: data = 6'b010101;
12'b11100011111001: data = 6'b000000;
12'b11100011111010: data = 6'b000000;
12'b11100011111011: data = 6'b000000;
12'b11100011111100: data = 6'b000000;
12'b11100011111101: data = 6'b000000;
12'b11100011111110: data = 6'b000000;
12'b11100011111111: data = 6'b000000;
12'b111000110000000: data = 6'b000000;
12'b111000110000001: data = 6'b000000;
12'b111000110000010: data = 6'b000000;
12'b111000110000011: data = 6'b000000;
12'b111000110000100: data = 6'b000000;
12'b111000110000101: data = 6'b000000;
12'b111000110000110: data = 6'b000000;
12'b111000110000111: data = 6'b000000;
12'b111000110001000: data = 6'b000000;
12'b111000110001001: data = 6'b000000;
12'b111000110001010: data = 6'b000000;
12'b111000110001011: data = 6'b000000;
12'b111000110001100: data = 6'b000000;
12'b111000110001101: data = 6'b000000;
12'b111000110001110: data = 6'b101010;
12'b111000110001111: data = 6'b101010;
12'b111000110010000: data = 6'b101010;
12'b111000110010001: data = 6'b101010;
12'b111000110010010: data = 6'b010101;
12'b111000110010011: data = 6'b010101;
12'b111000110010100: data = 6'b010101;
12'b111000110010101: data = 6'b010101;
12'b111000110010110: data = 6'b010101;
12'b111000110010111: data = 6'b010101;
12'b111000110011000: data = 6'b010101;
12'b111000110011001: data = 6'b010101;
12'b111000110011010: data = 6'b010101;
12'b111000110011011: data = 6'b010101;
12'b111000110011100: data = 6'b010101;
12'b111000110011101: data = 6'b010101;
12'b111000110011110: data = 6'b010101;
12'b111000110011111: data = 6'b010101;
12'b111000110100000: data = 6'b010101;
12'b111000110100001: data = 6'b010101;
12'b111000110100010: data = 6'b010101;
12'b111000110100011: data = 6'b010101;
12'b111000110100100: data = 6'b010101;
12'b111000110100101: data = 6'b010101;
12'b111000110100110: data = 6'b010101;
12'b111000110100111: data = 6'b010101;
12'b111000110101000: data = 6'b010101;
12'b111000110101001: data = 6'b010101;
12'b111000110101010: data = 6'b010101;
12'b1110010000000: data = 6'b010101;
12'b1110010000001: data = 6'b010101;
12'b1110010000010: data = 6'b010101;
12'b1110010000011: data = 6'b010101;
12'b1110010000100: data = 6'b010101;
12'b1110010000101: data = 6'b010101;
12'b1110010000110: data = 6'b010101;
12'b1110010000111: data = 6'b010101;
12'b1110010001000: data = 6'b010101;
12'b1110010001001: data = 6'b010101;
12'b1110010001010: data = 6'b010101;
12'b1110010001011: data = 6'b010101;
12'b1110010001100: data = 6'b010101;
12'b1110010001101: data = 6'b010101;
12'b1110010001110: data = 6'b010101;
12'b1110010001111: data = 6'b010101;
12'b1110010010000: data = 6'b010101;
12'b1110010010001: data = 6'b010101;
12'b1110010010010: data = 6'b010101;
12'b1110010010011: data = 6'b010101;
12'b1110010010100: data = 6'b010101;
12'b1110010010101: data = 6'b010101;
12'b1110010010110: data = 6'b010101;
12'b1110010010111: data = 6'b010101;
12'b1110010011000: data = 6'b010101;
12'b1110010011001: data = 6'b101010;
12'b1110010011010: data = 6'b101010;
12'b1110010011011: data = 6'b101010;
12'b1110010011100: data = 6'b010101;
12'b1110010011101: data = 6'b000000;
12'b1110010011110: data = 6'b000000;
12'b1110010011111: data = 6'b000000;
12'b1110010100000: data = 6'b000000;
12'b1110010100001: data = 6'b000000;
12'b1110010100010: data = 6'b000000;
12'b1110010100011: data = 6'b000000;
12'b1110010100100: data = 6'b000000;
12'b1110010100101: data = 6'b000000;
12'b1110010100110: data = 6'b000000;
12'b1110010100111: data = 6'b000000;
12'b1110010101000: data = 6'b000000;
12'b1110010101001: data = 6'b000000;
12'b1110010101010: data = 6'b000000;
12'b1110010101011: data = 6'b000000;
12'b1110010101100: data = 6'b000000;
12'b1110010101101: data = 6'b000000;
12'b1110010101110: data = 6'b000000;
12'b1110010101111: data = 6'b000000;
12'b1110010110000: data = 6'b000000;
12'b1110010110001: data = 6'b000000;
12'b1110010110010: data = 6'b000000;
12'b1110010110011: data = 6'b000000;
12'b1110010110100: data = 6'b000000;
12'b1110010110101: data = 6'b010101;
12'b1110010110110: data = 6'b010101;
12'b1110010110111: data = 6'b010101;
12'b1110010111000: data = 6'b010101;
12'b1110010111001: data = 6'b010101;
12'b1110010111010: data = 6'b010101;
12'b1110010111011: data = 6'b010101;
12'b1110010111100: data = 6'b010101;
12'b1110010111101: data = 6'b010101;
12'b1110010111110: data = 6'b010101;
12'b1110010111111: data = 6'b010101;
12'b11100101000000: data = 6'b010101;
12'b11100101000001: data = 6'b010101;
12'b11100101000010: data = 6'b010101;
12'b11100101000011: data = 6'b010101;
12'b11100101000100: data = 6'b010101;
12'b11100101000101: data = 6'b010101;
12'b11100101000110: data = 6'b010101;
12'b11100101000111: data = 6'b010101;
12'b11100101001000: data = 6'b010101;
12'b11100101001001: data = 6'b010101;
12'b11100101001010: data = 6'b010101;
12'b11100101001011: data = 6'b010101;
12'b11100101001100: data = 6'b010101;
12'b11100101001101: data = 6'b010101;
12'b11100101001110: data = 6'b010101;
12'b11100101001111: data = 6'b010101;
12'b11100101010000: data = 6'b010101;
12'b11100101010001: data = 6'b010101;
12'b11100101010010: data = 6'b010101;
12'b11100101010011: data = 6'b010101;
12'b11100101010100: data = 6'b010101;
12'b11100101010101: data = 6'b010101;
12'b11100101010110: data = 6'b010101;
12'b11100101010111: data = 6'b010101;
12'b11100101011000: data = 6'b010101;
12'b11100101011001: data = 6'b010101;
12'b11100101011010: data = 6'b010101;
12'b11100101011011: data = 6'b010101;
12'b11100101011100: data = 6'b010101;
12'b11100101011101: data = 6'b010101;
12'b11100101011110: data = 6'b010101;
12'b11100101011111: data = 6'b010101;
12'b11100101100000: data = 6'b010101;
12'b11100101100001: data = 6'b010101;
12'b11100101100010: data = 6'b010101;
12'b11100101100011: data = 6'b010101;
12'b11100101100100: data = 6'b010101;
12'b11100101100101: data = 6'b010101;
12'b11100101100110: data = 6'b010101;
12'b11100101100111: data = 6'b010101;
12'b11100101101000: data = 6'b010101;
12'b11100101101001: data = 6'b010101;
12'b11100101101010: data = 6'b010101;
12'b11100101101011: data = 6'b010101;
12'b11100101101100: data = 6'b010101;
12'b11100101101101: data = 6'b010101;
12'b11100101101110: data = 6'b010101;
12'b11100101101111: data = 6'b010101;
12'b11100101110000: data = 6'b010101;
12'b11100101110001: data = 6'b010101;
12'b11100101110010: data = 6'b010101;
12'b11100101110011: data = 6'b010101;
12'b11100101110100: data = 6'b010101;
12'b11100101110101: data = 6'b010101;
12'b11100101110110: data = 6'b010101;
12'b11100101110111: data = 6'b010101;
12'b11100101111000: data = 6'b000000;
12'b11100101111001: data = 6'b000000;
12'b11100101111010: data = 6'b010101;
12'b11100101111011: data = 6'b000000;
12'b11100101111100: data = 6'b000000;
12'b11100101111101: data = 6'b000000;
12'b11100101111110: data = 6'b000000;
12'b11100101111111: data = 6'b000000;
12'b111001010000000: data = 6'b000000;
12'b111001010000001: data = 6'b000000;
12'b111001010000010: data = 6'b000000;
12'b111001010000011: data = 6'b000000;
12'b111001010000100: data = 6'b000000;
12'b111001010000101: data = 6'b000000;
12'b111001010000110: data = 6'b000000;
12'b111001010000111: data = 6'b000000;
12'b111001010001000: data = 6'b000000;
12'b111001010001001: data = 6'b000000;
12'b111001010001010: data = 6'b000000;
12'b111001010001011: data = 6'b000000;
12'b111001010001100: data = 6'b000000;
12'b111001010001101: data = 6'b000000;
12'b111001010001110: data = 6'b101010;
12'b111001010001111: data = 6'b101010;
12'b111001010010000: data = 6'b101010;
12'b111001010010001: data = 6'b101010;
12'b111001010010010: data = 6'b010101;
12'b111001010010011: data = 6'b010101;
12'b111001010010100: data = 6'b010101;
12'b111001010010101: data = 6'b010101;
12'b111001010010110: data = 6'b010101;
12'b111001010010111: data = 6'b010101;
12'b111001010011000: data = 6'b010101;
12'b111001010011001: data = 6'b010101;
12'b111001010011010: data = 6'b010101;
12'b111001010011011: data = 6'b010101;
12'b111001010011100: data = 6'b010101;
12'b111001010011101: data = 6'b010101;
12'b111001010011110: data = 6'b010101;
12'b111001010011111: data = 6'b010101;
12'b111001010100000: data = 6'b010101;
12'b111001010100001: data = 6'b010101;
12'b111001010100010: data = 6'b010101;
12'b111001010100011: data = 6'b010101;
12'b111001010100100: data = 6'b010101;
12'b111001010100101: data = 6'b010101;
12'b111001010100110: data = 6'b010101;
12'b111001010100111: data = 6'b010101;
12'b111001010101000: data = 6'b010101;
12'b111001010101001: data = 6'b010101;
12'b111001010101010: data = 6'b010101;
12'b1110011000000: data = 6'b010101;
12'b1110011000001: data = 6'b010101;
12'b1110011000010: data = 6'b010101;
12'b1110011000011: data = 6'b010101;
12'b1110011000100: data = 6'b010101;
12'b1110011000101: data = 6'b010101;
12'b1110011000110: data = 6'b010101;
12'b1110011000111: data = 6'b010101;
12'b1110011001000: data = 6'b010101;
12'b1110011001001: data = 6'b010101;
12'b1110011001010: data = 6'b010101;
12'b1110011001011: data = 6'b010101;
12'b1110011001100: data = 6'b010101;
12'b1110011001101: data = 6'b010101;
12'b1110011001110: data = 6'b010101;
12'b1110011001111: data = 6'b010101;
12'b1110011010000: data = 6'b010101;
12'b1110011010001: data = 6'b010101;
12'b1110011010010: data = 6'b010101;
12'b1110011010011: data = 6'b010101;
12'b1110011010100: data = 6'b010101;
12'b1110011010101: data = 6'b010101;
12'b1110011010110: data = 6'b010101;
12'b1110011010111: data = 6'b010101;
12'b1110011011000: data = 6'b010101;
12'b1110011011001: data = 6'b101010;
12'b1110011011010: data = 6'b101010;
12'b1110011011011: data = 6'b101010;
12'b1110011011100: data = 6'b010101;
12'b1110011011101: data = 6'b000000;
12'b1110011011110: data = 6'b000000;
12'b1110011011111: data = 6'b000000;
12'b1110011100000: data = 6'b000000;
12'b1110011100001: data = 6'b000000;
12'b1110011100010: data = 6'b000000;
12'b1110011100011: data = 6'b000000;
12'b1110011100100: data = 6'b000000;
12'b1110011100101: data = 6'b000000;
12'b1110011100110: data = 6'b000000;
12'b1110011100111: data = 6'b000000;
12'b1110011101000: data = 6'b000000;
12'b1110011101001: data = 6'b000000;
12'b1110011101010: data = 6'b000000;
12'b1110011101011: data = 6'b000000;
12'b1110011101100: data = 6'b000000;
12'b1110011101101: data = 6'b000000;
12'b1110011101110: data = 6'b000000;
12'b1110011101111: data = 6'b000000;
12'b1110011110000: data = 6'b000000;
12'b1110011110001: data = 6'b000000;
12'b1110011110010: data = 6'b000000;
12'b1110011110011: data = 6'b000000;
12'b1110011110100: data = 6'b000000;
12'b1110011110101: data = 6'b010101;
12'b1110011110110: data = 6'b000000;
12'b1110011110111: data = 6'b010101;
12'b1110011111000: data = 6'b010101;
12'b1110011111001: data = 6'b010101;
12'b1110011111010: data = 6'b010101;
12'b1110011111011: data = 6'b010101;
12'b1110011111100: data = 6'b010101;
12'b1110011111101: data = 6'b010101;
12'b1110011111110: data = 6'b010101;
12'b1110011111111: data = 6'b010101;
12'b11100111000000: data = 6'b010101;
12'b11100111000001: data = 6'b010101;
12'b11100111000010: data = 6'b010101;
12'b11100111000011: data = 6'b010101;
12'b11100111000100: data = 6'b010101;
12'b11100111000101: data = 6'b010101;
12'b11100111000110: data = 6'b010101;
12'b11100111000111: data = 6'b010101;
12'b11100111001000: data = 6'b010101;
12'b11100111001001: data = 6'b010101;
12'b11100111001010: data = 6'b010101;
12'b11100111001011: data = 6'b010101;
12'b11100111001100: data = 6'b010101;
12'b11100111001101: data = 6'b010101;
12'b11100111001110: data = 6'b010101;
12'b11100111001111: data = 6'b010101;
12'b11100111010000: data = 6'b010101;
12'b11100111010001: data = 6'b010101;
12'b11100111010010: data = 6'b010101;
12'b11100111010011: data = 6'b010101;
12'b11100111010100: data = 6'b010101;
12'b11100111010101: data = 6'b010101;
12'b11100111010110: data = 6'b010101;
12'b11100111010111: data = 6'b010101;
12'b11100111011000: data = 6'b010101;
12'b11100111011001: data = 6'b010101;
12'b11100111011010: data = 6'b010101;
12'b11100111011011: data = 6'b010101;
12'b11100111011100: data = 6'b010101;
12'b11100111011101: data = 6'b010101;
12'b11100111011110: data = 6'b010101;
12'b11100111011111: data = 6'b010101;
12'b11100111100000: data = 6'b010101;
12'b11100111100001: data = 6'b010101;
12'b11100111100010: data = 6'b010101;
12'b11100111100011: data = 6'b010101;
12'b11100111100100: data = 6'b010101;
12'b11100111100101: data = 6'b010101;
12'b11100111100110: data = 6'b010101;
12'b11100111100111: data = 6'b010101;
12'b11100111101000: data = 6'b010101;
12'b11100111101001: data = 6'b010101;
12'b11100111101010: data = 6'b010101;
12'b11100111101011: data = 6'b010101;
12'b11100111101100: data = 6'b010101;
12'b11100111101101: data = 6'b010101;
12'b11100111101110: data = 6'b010101;
12'b11100111101111: data = 6'b010101;
12'b11100111110000: data = 6'b010101;
12'b11100111110001: data = 6'b010101;
12'b11100111110010: data = 6'b010101;
12'b11100111110011: data = 6'b010101;
12'b11100111110100: data = 6'b010101;
12'b11100111110101: data = 6'b010101;
12'b11100111110110: data = 6'b010101;
12'b11100111110111: data = 6'b010101;
12'b11100111111000: data = 6'b010101;
12'b11100111111001: data = 6'b000000;
12'b11100111111010: data = 6'b000000;
12'b11100111111011: data = 6'b000000;
12'b11100111111100: data = 6'b000000;
12'b11100111111101: data = 6'b000000;
12'b11100111111110: data = 6'b000000;
12'b11100111111111: data = 6'b000000;
12'b111001110000000: data = 6'b000000;
12'b111001110000001: data = 6'b000000;
12'b111001110000010: data = 6'b000000;
12'b111001110000011: data = 6'b000000;
12'b111001110000100: data = 6'b000000;
12'b111001110000101: data = 6'b000000;
12'b111001110000110: data = 6'b000000;
12'b111001110000111: data = 6'b000000;
12'b111001110001000: data = 6'b000000;
12'b111001110001001: data = 6'b000000;
12'b111001110001010: data = 6'b000000;
12'b111001110001011: data = 6'b000000;
12'b111001110001100: data = 6'b000000;
12'b111001110001101: data = 6'b000000;
12'b111001110001110: data = 6'b101010;
12'b111001110001111: data = 6'b101010;
12'b111001110010000: data = 6'b101010;
12'b111001110010001: data = 6'b101010;
12'b111001110010010: data = 6'b010101;
12'b111001110010011: data = 6'b010101;
12'b111001110010100: data = 6'b010101;
12'b111001110010101: data = 6'b010101;
12'b111001110010110: data = 6'b010101;
12'b111001110010111: data = 6'b010101;
12'b111001110011000: data = 6'b010101;
12'b111001110011001: data = 6'b010101;
12'b111001110011010: data = 6'b010101;
12'b111001110011011: data = 6'b010101;
12'b111001110011100: data = 6'b010101;
12'b111001110011101: data = 6'b010101;
12'b111001110011110: data = 6'b010101;
12'b111001110011111: data = 6'b010101;
12'b111001110100000: data = 6'b010101;
12'b111001110100001: data = 6'b010101;
12'b111001110100010: data = 6'b010101;
12'b111001110100011: data = 6'b010101;
12'b111001110100100: data = 6'b010101;
12'b111001110100101: data = 6'b010101;
12'b111001110100110: data = 6'b010101;
12'b111001110100111: data = 6'b010101;
12'b111001110101000: data = 6'b010101;
12'b111001110101001: data = 6'b010101;
12'b111001110101010: data = 6'b010101;
12'b1110100000000: data = 6'b010101;
12'b1110100000001: data = 6'b010101;
12'b1110100000010: data = 6'b010101;
12'b1110100000011: data = 6'b010101;
12'b1110100000100: data = 6'b010101;
12'b1110100000101: data = 6'b010101;
12'b1110100000110: data = 6'b010101;
12'b1110100000111: data = 6'b010101;
12'b1110100001000: data = 6'b010101;
12'b1110100001001: data = 6'b010101;
12'b1110100001010: data = 6'b010101;
12'b1110100001011: data = 6'b010101;
12'b1110100001100: data = 6'b010101;
12'b1110100001101: data = 6'b010101;
12'b1110100001110: data = 6'b010101;
12'b1110100001111: data = 6'b010101;
12'b1110100010000: data = 6'b010101;
12'b1110100010001: data = 6'b010101;
12'b1110100010010: data = 6'b010101;
12'b1110100010011: data = 6'b010101;
12'b1110100010100: data = 6'b010101;
12'b1110100010101: data = 6'b010101;
12'b1110100010110: data = 6'b010101;
12'b1110100010111: data = 6'b010101;
12'b1110100011000: data = 6'b010101;
12'b1110100011001: data = 6'b101010;
12'b1110100011010: data = 6'b101010;
12'b1110100011011: data = 6'b101010;
12'b1110100011100: data = 6'b010101;
12'b1110100011101: data = 6'b000000;
12'b1110100011110: data = 6'b000000;
12'b1110100011111: data = 6'b000000;
12'b1110100100000: data = 6'b000000;
12'b1110100100001: data = 6'b000000;
12'b1110100100010: data = 6'b000000;
12'b1110100100011: data = 6'b000000;
12'b1110100100100: data = 6'b000000;
12'b1110100100101: data = 6'b000000;
12'b1110100100110: data = 6'b000000;
12'b1110100100111: data = 6'b000000;
12'b1110100101000: data = 6'b000000;
12'b1110100101001: data = 6'b000000;
12'b1110100101010: data = 6'b000000;
12'b1110100101011: data = 6'b000000;
12'b1110100101100: data = 6'b000000;
12'b1110100101101: data = 6'b000000;
12'b1110100101110: data = 6'b000000;
12'b1110100101111: data = 6'b000000;
12'b1110100110000: data = 6'b000000;
12'b1110100110001: data = 6'b000000;
12'b1110100110010: data = 6'b000000;
12'b1110100110011: data = 6'b000000;
12'b1110100110100: data = 6'b000000;
12'b1110100110101: data = 6'b010101;
12'b1110100110110: data = 6'b010101;
12'b1110100110111: data = 6'b010101;
12'b1110100111000: data = 6'b010101;
12'b1110100111001: data = 6'b010101;
12'b1110100111010: data = 6'b010101;
12'b1110100111011: data = 6'b010101;
12'b1110100111100: data = 6'b010101;
12'b1110100111101: data = 6'b010101;
12'b1110100111110: data = 6'b010101;
12'b1110100111111: data = 6'b010101;
12'b11101001000000: data = 6'b010101;
12'b11101001000001: data = 6'b010101;
12'b11101001000010: data = 6'b010101;
12'b11101001000011: data = 6'b010101;
12'b11101001000100: data = 6'b010101;
12'b11101001000101: data = 6'b010101;
12'b11101001000110: data = 6'b010101;
12'b11101001000111: data = 6'b010101;
12'b11101001001000: data = 6'b010101;
12'b11101001001001: data = 6'b010101;
12'b11101001001010: data = 6'b010101;
12'b11101001001011: data = 6'b010101;
12'b11101001001100: data = 6'b010101;
12'b11101001001101: data = 6'b010101;
12'b11101001001110: data = 6'b010101;
12'b11101001001111: data = 6'b010101;
12'b11101001010000: data = 6'b010101;
12'b11101001010001: data = 6'b010101;
12'b11101001010010: data = 6'b010101;
12'b11101001010011: data = 6'b010101;
12'b11101001010100: data = 6'b010101;
12'b11101001010101: data = 6'b010101;
12'b11101001010110: data = 6'b010101;
12'b11101001010111: data = 6'b010101;
12'b11101001011000: data = 6'b010101;
12'b11101001011001: data = 6'b010101;
12'b11101001011010: data = 6'b010101;
12'b11101001011011: data = 6'b010101;
12'b11101001011100: data = 6'b010101;
12'b11101001011101: data = 6'b010101;
12'b11101001011110: data = 6'b010101;
12'b11101001011111: data = 6'b010101;
12'b11101001100000: data = 6'b010101;
12'b11101001100001: data = 6'b010101;
12'b11101001100010: data = 6'b010101;
12'b11101001100011: data = 6'b010101;
12'b11101001100100: data = 6'b010101;
12'b11101001100101: data = 6'b010101;
12'b11101001100110: data = 6'b010101;
12'b11101001100111: data = 6'b010101;
12'b11101001101000: data = 6'b010101;
12'b11101001101001: data = 6'b010101;
12'b11101001101010: data = 6'b010101;
12'b11101001101011: data = 6'b010101;
12'b11101001101100: data = 6'b010101;
12'b11101001101101: data = 6'b010101;
12'b11101001101110: data = 6'b010101;
12'b11101001101111: data = 6'b010101;
12'b11101001110000: data = 6'b010101;
12'b11101001110001: data = 6'b010101;
12'b11101001110010: data = 6'b010101;
12'b11101001110011: data = 6'b010101;
12'b11101001110100: data = 6'b010101;
12'b11101001110101: data = 6'b010101;
12'b11101001110110: data = 6'b010101;
12'b11101001110111: data = 6'b010101;
12'b11101001111000: data = 6'b000000;
12'b11101001111001: data = 6'b010101;
12'b11101001111010: data = 6'b000000;
12'b11101001111011: data = 6'b000000;
12'b11101001111100: data = 6'b000000;
12'b11101001111101: data = 6'b000000;
12'b11101001111110: data = 6'b000000;
12'b11101001111111: data = 6'b000000;
12'b111010010000000: data = 6'b000000;
12'b111010010000001: data = 6'b000000;
12'b111010010000010: data = 6'b000000;
12'b111010010000011: data = 6'b000000;
12'b111010010000100: data = 6'b000000;
12'b111010010000101: data = 6'b000000;
12'b111010010000110: data = 6'b000000;
12'b111010010000111: data = 6'b000000;
12'b111010010001000: data = 6'b000000;
12'b111010010001001: data = 6'b000000;
12'b111010010001010: data = 6'b000000;
12'b111010010001011: data = 6'b000000;
12'b111010010001100: data = 6'b000000;
12'b111010010001101: data = 6'b000000;
12'b111010010001110: data = 6'b101010;
12'b111010010001111: data = 6'b101010;
12'b111010010010000: data = 6'b101010;
12'b111010010010001: data = 6'b101010;
12'b111010010010010: data = 6'b010101;
12'b111010010010011: data = 6'b010101;
12'b111010010010100: data = 6'b010101;
12'b111010010010101: data = 6'b010101;
12'b111010010010110: data = 6'b010101;
12'b111010010010111: data = 6'b010101;
12'b111010010011000: data = 6'b010101;
12'b111010010011001: data = 6'b010101;
12'b111010010011010: data = 6'b010101;
12'b111010010011011: data = 6'b010101;
12'b111010010011100: data = 6'b010101;
12'b111010010011101: data = 6'b010101;
12'b111010010011110: data = 6'b010101;
12'b111010010011111: data = 6'b010101;
12'b111010010100000: data = 6'b010101;
12'b111010010100001: data = 6'b010101;
12'b111010010100010: data = 6'b010101;
12'b111010010100011: data = 6'b010101;
12'b111010010100100: data = 6'b010101;
12'b111010010100101: data = 6'b010101;
12'b111010010100110: data = 6'b010101;
12'b111010010100111: data = 6'b010101;
12'b111010010101000: data = 6'b010101;
12'b111010010101001: data = 6'b010101;
12'b111010010101010: data = 6'b010101;
12'b1110101000000: data = 6'b010101;
12'b1110101000001: data = 6'b010101;
12'b1110101000010: data = 6'b010101;
12'b1110101000011: data = 6'b010101;
12'b1110101000100: data = 6'b010101;
12'b1110101000101: data = 6'b010101;
12'b1110101000110: data = 6'b010101;
12'b1110101000111: data = 6'b010101;
12'b1110101001000: data = 6'b010101;
12'b1110101001001: data = 6'b010101;
12'b1110101001010: data = 6'b010101;
12'b1110101001011: data = 6'b010101;
12'b1110101001100: data = 6'b010101;
12'b1110101001101: data = 6'b010101;
12'b1110101001110: data = 6'b010101;
12'b1110101001111: data = 6'b010101;
12'b1110101010000: data = 6'b010101;
12'b1110101010001: data = 6'b010101;
12'b1110101010010: data = 6'b010101;
12'b1110101010011: data = 6'b010101;
12'b1110101010100: data = 6'b010101;
12'b1110101010101: data = 6'b010101;
12'b1110101010110: data = 6'b010101;
12'b1110101010111: data = 6'b010101;
12'b1110101011000: data = 6'b010101;
12'b1110101011001: data = 6'b101010;
12'b1110101011010: data = 6'b101010;
12'b1110101011011: data = 6'b101010;
12'b1110101011100: data = 6'b010101;
12'b1110101011101: data = 6'b000000;
12'b1110101011110: data = 6'b000000;
12'b1110101011111: data = 6'b000000;
12'b1110101100000: data = 6'b000000;
12'b1110101100001: data = 6'b000000;
12'b1110101100010: data = 6'b000000;
12'b1110101100011: data = 6'b000000;
12'b1110101100100: data = 6'b000000;
12'b1110101100101: data = 6'b000000;
12'b1110101100110: data = 6'b000000;
12'b1110101100111: data = 6'b000000;
12'b1110101101000: data = 6'b000000;
12'b1110101101001: data = 6'b000000;
12'b1110101101010: data = 6'b000000;
12'b1110101101011: data = 6'b000000;
12'b1110101101100: data = 6'b000000;
12'b1110101101101: data = 6'b000000;
12'b1110101101110: data = 6'b000000;
12'b1110101101111: data = 6'b000000;
12'b1110101110000: data = 6'b000000;
12'b1110101110001: data = 6'b000000;
12'b1110101110010: data = 6'b000000;
12'b1110101110011: data = 6'b000000;
12'b1110101110100: data = 6'b000000;
12'b1110101110101: data = 6'b000000;
12'b1110101110110: data = 6'b010101;
12'b1110101110111: data = 6'b010101;
12'b1110101111000: data = 6'b010101;
12'b1110101111001: data = 6'b010101;
12'b1110101111010: data = 6'b010101;
12'b1110101111011: data = 6'b010101;
12'b1110101111100: data = 6'b010101;
12'b1110101111101: data = 6'b010101;
12'b1110101111110: data = 6'b010101;
12'b1110101111111: data = 6'b010101;
12'b11101011000000: data = 6'b010101;
12'b11101011000001: data = 6'b010101;
12'b11101011000010: data = 6'b010101;
12'b11101011000011: data = 6'b010101;
12'b11101011000100: data = 6'b010101;
12'b11101011000101: data = 6'b010101;
12'b11101011000110: data = 6'b010101;
12'b11101011000111: data = 6'b010101;
12'b11101011001000: data = 6'b010101;
12'b11101011001001: data = 6'b010101;
12'b11101011001010: data = 6'b010101;
12'b11101011001011: data = 6'b010101;
12'b11101011001100: data = 6'b010101;
12'b11101011001101: data = 6'b010101;
12'b11101011001110: data = 6'b010101;
12'b11101011001111: data = 6'b010101;
12'b11101011010000: data = 6'b010101;
12'b11101011010001: data = 6'b010101;
12'b11101011010010: data = 6'b010101;
12'b11101011010011: data = 6'b010101;
12'b11101011010100: data = 6'b010101;
12'b11101011010101: data = 6'b010101;
12'b11101011010110: data = 6'b010101;
12'b11101011010111: data = 6'b010101;
12'b11101011011000: data = 6'b010101;
12'b11101011011001: data = 6'b010101;
12'b11101011011010: data = 6'b010101;
12'b11101011011011: data = 6'b010101;
12'b11101011011100: data = 6'b010101;
12'b11101011011101: data = 6'b010101;
12'b11101011011110: data = 6'b010101;
12'b11101011011111: data = 6'b010101;
12'b11101011100000: data = 6'b010101;
12'b11101011100001: data = 6'b010101;
12'b11101011100010: data = 6'b010101;
12'b11101011100011: data = 6'b010101;
12'b11101011100100: data = 6'b010101;
12'b11101011100101: data = 6'b010101;
12'b11101011100110: data = 6'b010101;
12'b11101011100111: data = 6'b010101;
12'b11101011101000: data = 6'b010101;
12'b11101011101001: data = 6'b010101;
12'b11101011101010: data = 6'b010101;
12'b11101011101011: data = 6'b010101;
12'b11101011101100: data = 6'b010101;
12'b11101011101101: data = 6'b010101;
12'b11101011101110: data = 6'b010101;
12'b11101011101111: data = 6'b010101;
12'b11101011110000: data = 6'b010101;
12'b11101011110001: data = 6'b010101;
12'b11101011110010: data = 6'b010101;
12'b11101011110011: data = 6'b010101;
12'b11101011110100: data = 6'b010101;
12'b11101011110101: data = 6'b010101;
12'b11101011110110: data = 6'b010101;
12'b11101011110111: data = 6'b010101;
12'b11101011111000: data = 6'b010101;
12'b11101011111001: data = 6'b000000;
12'b11101011111010: data = 6'b000000;
12'b11101011111011: data = 6'b000000;
12'b11101011111100: data = 6'b000000;
12'b11101011111101: data = 6'b000000;
12'b11101011111110: data = 6'b000000;
12'b11101011111111: data = 6'b000000;
12'b111010110000000: data = 6'b000000;
12'b111010110000001: data = 6'b000000;
12'b111010110000010: data = 6'b000000;
12'b111010110000011: data = 6'b000000;
12'b111010110000100: data = 6'b000000;
12'b111010110000101: data = 6'b000000;
12'b111010110000110: data = 6'b000000;
12'b111010110000111: data = 6'b000000;
12'b111010110001000: data = 6'b000000;
12'b111010110001001: data = 6'b000000;
12'b111010110001010: data = 6'b000000;
12'b111010110001011: data = 6'b000000;
12'b111010110001100: data = 6'b000000;
12'b111010110001101: data = 6'b000000;
12'b111010110001110: data = 6'b101010;
12'b111010110001111: data = 6'b101010;
12'b111010110010000: data = 6'b101010;
12'b111010110010001: data = 6'b101010;
12'b111010110010010: data = 6'b010101;
12'b111010110010011: data = 6'b010101;
12'b111010110010100: data = 6'b010101;
12'b111010110010101: data = 6'b010101;
12'b111010110010110: data = 6'b010101;
12'b111010110010111: data = 6'b010101;
12'b111010110011000: data = 6'b010101;
12'b111010110011001: data = 6'b010101;
12'b111010110011010: data = 6'b010101;
12'b111010110011011: data = 6'b010101;
12'b111010110011100: data = 6'b010101;
12'b111010110011101: data = 6'b010101;
12'b111010110011110: data = 6'b010101;
12'b111010110011111: data = 6'b010101;
12'b111010110100000: data = 6'b010101;
12'b111010110100001: data = 6'b010101;
12'b111010110100010: data = 6'b010101;
12'b111010110100011: data = 6'b010101;
12'b111010110100100: data = 6'b010101;
12'b111010110100101: data = 6'b010101;
12'b111010110100110: data = 6'b010101;
12'b111010110100111: data = 6'b010101;
12'b111010110101000: data = 6'b010101;
12'b111010110101001: data = 6'b010101;
12'b111010110101010: data = 6'b010101;
12'b1110110000000: data = 6'b010101;
12'b1110110000001: data = 6'b010101;
12'b1110110000010: data = 6'b010101;
12'b1110110000011: data = 6'b010101;
12'b1110110000100: data = 6'b010101;
12'b1110110000101: data = 6'b010101;
12'b1110110000110: data = 6'b010101;
12'b1110110000111: data = 6'b010101;
12'b1110110001000: data = 6'b010101;
12'b1110110001001: data = 6'b010101;
12'b1110110001010: data = 6'b010101;
12'b1110110001011: data = 6'b010101;
12'b1110110001100: data = 6'b010101;
12'b1110110001101: data = 6'b010101;
12'b1110110001110: data = 6'b010101;
12'b1110110001111: data = 6'b010101;
12'b1110110010000: data = 6'b010101;
12'b1110110010001: data = 6'b010101;
12'b1110110010010: data = 6'b010101;
12'b1110110010011: data = 6'b010101;
12'b1110110010100: data = 6'b010101;
12'b1110110010101: data = 6'b010101;
12'b1110110010110: data = 6'b010101;
12'b1110110010111: data = 6'b010101;
12'b1110110011000: data = 6'b010101;
12'b1110110011001: data = 6'b101010;
12'b1110110011010: data = 6'b101010;
12'b1110110011011: data = 6'b101010;
12'b1110110011100: data = 6'b010101;
12'b1110110011101: data = 6'b000000;
12'b1110110011110: data = 6'b000000;
12'b1110110011111: data = 6'b000000;
12'b1110110100000: data = 6'b000000;
12'b1110110100001: data = 6'b000000;
12'b1110110100010: data = 6'b000000;
12'b1110110100011: data = 6'b000000;
12'b1110110100100: data = 6'b000000;
12'b1110110100101: data = 6'b000000;
12'b1110110100110: data = 6'b000000;
12'b1110110100111: data = 6'b000000;
12'b1110110101000: data = 6'b000000;
12'b1110110101001: data = 6'b000000;
12'b1110110101010: data = 6'b000000;
12'b1110110101011: data = 6'b000000;
12'b1110110101100: data = 6'b000000;
12'b1110110101101: data = 6'b000000;
12'b1110110101110: data = 6'b000000;
12'b1110110101111: data = 6'b000000;
12'b1110110110000: data = 6'b000000;
12'b1110110110001: data = 6'b000000;
12'b1110110110010: data = 6'b000000;
12'b1110110110011: data = 6'b000000;
12'b1110110110100: data = 6'b000000;
12'b1110110110101: data = 6'b010101;
12'b1110110110110: data = 6'b010101;
12'b1110110110111: data = 6'b010101;
12'b1110110111000: data = 6'b010101;
12'b1110110111001: data = 6'b010101;
12'b1110110111010: data = 6'b010101;
12'b1110110111011: data = 6'b010101;
12'b1110110111100: data = 6'b010101;
12'b1110110111101: data = 6'b010101;
12'b1110110111110: data = 6'b010101;
12'b1110110111111: data = 6'b010101;
12'b11101101000000: data = 6'b010101;
12'b11101101000001: data = 6'b010101;
12'b11101101000010: data = 6'b010101;
12'b11101101000011: data = 6'b010101;
12'b11101101000100: data = 6'b010101;
12'b11101101000101: data = 6'b010101;
12'b11101101000110: data = 6'b010101;
12'b11101101000111: data = 6'b010101;
12'b11101101001000: data = 6'b010101;
12'b11101101001001: data = 6'b010101;
12'b11101101001010: data = 6'b010101;
12'b11101101001011: data = 6'b010101;
12'b11101101001100: data = 6'b010101;
12'b11101101001101: data = 6'b010101;
12'b11101101001110: data = 6'b010101;
12'b11101101001111: data = 6'b010101;
12'b11101101010000: data = 6'b010101;
12'b11101101010001: data = 6'b010101;
12'b11101101010010: data = 6'b010101;
12'b11101101010011: data = 6'b010101;
12'b11101101010100: data = 6'b010101;
12'b11101101010101: data = 6'b010101;
12'b11101101010110: data = 6'b010101;
12'b11101101010111: data = 6'b010101;
12'b11101101011000: data = 6'b010101;
12'b11101101011001: data = 6'b010101;
12'b11101101011010: data = 6'b010101;
12'b11101101011011: data = 6'b010101;
12'b11101101011100: data = 6'b010101;
12'b11101101011101: data = 6'b010101;
12'b11101101011110: data = 6'b010101;
12'b11101101011111: data = 6'b010101;
12'b11101101100000: data = 6'b010101;
12'b11101101100001: data = 6'b010101;
12'b11101101100010: data = 6'b010101;
12'b11101101100011: data = 6'b010101;
12'b11101101100100: data = 6'b010101;
12'b11101101100101: data = 6'b010101;
12'b11101101100110: data = 6'b010101;
12'b11101101100111: data = 6'b010101;
12'b11101101101000: data = 6'b010101;
12'b11101101101001: data = 6'b010101;
12'b11101101101010: data = 6'b010101;
12'b11101101101011: data = 6'b010101;
12'b11101101101100: data = 6'b010101;
12'b11101101101101: data = 6'b010101;
12'b11101101101110: data = 6'b010101;
12'b11101101101111: data = 6'b010101;
12'b11101101110000: data = 6'b010101;
12'b11101101110001: data = 6'b010101;
12'b11101101110010: data = 6'b010101;
12'b11101101110011: data = 6'b010101;
12'b11101101110100: data = 6'b010101;
12'b11101101110101: data = 6'b010101;
12'b11101101110110: data = 6'b010101;
12'b11101101110111: data = 6'b000000;
12'b11101101111000: data = 6'b010101;
12'b11101101111001: data = 6'b000000;
12'b11101101111010: data = 6'b000000;
12'b11101101111011: data = 6'b000000;
12'b11101101111100: data = 6'b000000;
12'b11101101111101: data = 6'b000000;
12'b11101101111110: data = 6'b000000;
12'b11101101111111: data = 6'b000000;
12'b111011010000000: data = 6'b000000;
12'b111011010000001: data = 6'b000000;
12'b111011010000010: data = 6'b000000;
12'b111011010000011: data = 6'b000000;
12'b111011010000100: data = 6'b000000;
12'b111011010000101: data = 6'b000000;
12'b111011010000110: data = 6'b000000;
12'b111011010000111: data = 6'b000000;
12'b111011010001000: data = 6'b000000;
12'b111011010001001: data = 6'b000000;
12'b111011010001010: data = 6'b000000;
12'b111011010001011: data = 6'b000000;
12'b111011010001100: data = 6'b000000;
12'b111011010001101: data = 6'b000000;
12'b111011010001110: data = 6'b101010;
12'b111011010001111: data = 6'b101010;
12'b111011010010000: data = 6'b101010;
12'b111011010010001: data = 6'b101010;
12'b111011010010010: data = 6'b010101;
12'b111011010010011: data = 6'b010101;
12'b111011010010100: data = 6'b010101;
12'b111011010010101: data = 6'b010101;
12'b111011010010110: data = 6'b010101;
12'b111011010010111: data = 6'b010101;
12'b111011010011000: data = 6'b010101;
12'b111011010011001: data = 6'b010101;
12'b111011010011010: data = 6'b010101;
12'b111011010011011: data = 6'b010101;
12'b111011010011100: data = 6'b010101;
12'b111011010011101: data = 6'b010101;
12'b111011010011110: data = 6'b010101;
12'b111011010011111: data = 6'b010101;
12'b111011010100000: data = 6'b010101;
12'b111011010100001: data = 6'b010101;
12'b111011010100010: data = 6'b010101;
12'b111011010100011: data = 6'b010101;
12'b111011010100100: data = 6'b010101;
12'b111011010100101: data = 6'b010101;
12'b111011010100110: data = 6'b010101;
12'b111011010100111: data = 6'b010101;
12'b111011010101000: data = 6'b010101;
12'b111011010101001: data = 6'b010101;
12'b111011010101010: data = 6'b010101;
12'b1110111000000: data = 6'b010101;
12'b1110111000001: data = 6'b010101;
12'b1110111000010: data = 6'b010101;
12'b1110111000011: data = 6'b010101;
12'b1110111000100: data = 6'b010101;
12'b1110111000101: data = 6'b010101;
12'b1110111000110: data = 6'b010101;
12'b1110111000111: data = 6'b010101;
12'b1110111001000: data = 6'b010101;
12'b1110111001001: data = 6'b010101;
12'b1110111001010: data = 6'b010101;
12'b1110111001011: data = 6'b010101;
12'b1110111001100: data = 6'b010101;
12'b1110111001101: data = 6'b010101;
12'b1110111001110: data = 6'b010101;
12'b1110111001111: data = 6'b010101;
12'b1110111010000: data = 6'b010101;
12'b1110111010001: data = 6'b010101;
12'b1110111010010: data = 6'b010101;
12'b1110111010011: data = 6'b010101;
12'b1110111010100: data = 6'b010101;
12'b1110111010101: data = 6'b010101;
12'b1110111010110: data = 6'b010101;
12'b1110111010111: data = 6'b010101;
12'b1110111011000: data = 6'b010101;
12'b1110111011001: data = 6'b101010;
12'b1110111011010: data = 6'b101010;
12'b1110111011011: data = 6'b101010;
12'b1110111011100: data = 6'b101001;
12'b1110111011101: data = 6'b000000;
12'b1110111011110: data = 6'b000000;
12'b1110111011111: data = 6'b000000;
12'b1110111100000: data = 6'b000000;
12'b1110111100001: data = 6'b000000;
12'b1110111100010: data = 6'b000000;
12'b1110111100011: data = 6'b000000;
12'b1110111100100: data = 6'b000000;
12'b1110111100101: data = 6'b000000;
12'b1110111100110: data = 6'b000000;
12'b1110111100111: data = 6'b000000;
12'b1110111101000: data = 6'b000000;
12'b1110111101001: data = 6'b000000;
12'b1110111101010: data = 6'b000000;
12'b1110111101011: data = 6'b000000;
12'b1110111101100: data = 6'b000000;
12'b1110111101101: data = 6'b000000;
12'b1110111101110: data = 6'b000000;
12'b1110111101111: data = 6'b000000;
12'b1110111110000: data = 6'b000000;
12'b1110111110001: data = 6'b000000;
12'b1110111110010: data = 6'b000000;
12'b1110111110011: data = 6'b000000;
12'b1110111110100: data = 6'b000000;
12'b1110111110101: data = 6'b010101;
12'b1110111110110: data = 6'b010101;
12'b1110111110111: data = 6'b010101;
12'b1110111111000: data = 6'b010101;
12'b1110111111001: data = 6'b010101;
12'b1110111111010: data = 6'b010101;
12'b1110111111011: data = 6'b010101;
12'b1110111111100: data = 6'b010101;
12'b1110111111101: data = 6'b010101;
12'b1110111111110: data = 6'b010101;
12'b1110111111111: data = 6'b010101;
12'b11101111000000: data = 6'b010101;
12'b11101111000001: data = 6'b010101;
12'b11101111000010: data = 6'b010101;
12'b11101111000011: data = 6'b010101;
12'b11101111000100: data = 6'b010101;
12'b11101111000101: data = 6'b010101;
12'b11101111000110: data = 6'b010101;
12'b11101111000111: data = 6'b010101;
12'b11101111001000: data = 6'b010101;
12'b11101111001001: data = 6'b010101;
12'b11101111001010: data = 6'b010101;
12'b11101111001011: data = 6'b010101;
12'b11101111001100: data = 6'b010101;
12'b11101111001101: data = 6'b010101;
12'b11101111001110: data = 6'b010101;
12'b11101111001111: data = 6'b010101;
12'b11101111010000: data = 6'b010101;
12'b11101111010001: data = 6'b010101;
12'b11101111010010: data = 6'b010101;
12'b11101111010011: data = 6'b010101;
12'b11101111010100: data = 6'b010101;
12'b11101111010101: data = 6'b010101;
12'b11101111010110: data = 6'b010101;
12'b11101111010111: data = 6'b010101;
12'b11101111011000: data = 6'b010101;
12'b11101111011001: data = 6'b010101;
12'b11101111011010: data = 6'b010101;
12'b11101111011011: data = 6'b010101;
12'b11101111011100: data = 6'b010101;
12'b11101111011101: data = 6'b010101;
12'b11101111011110: data = 6'b010101;
12'b11101111011111: data = 6'b010101;
12'b11101111100000: data = 6'b010101;
12'b11101111100001: data = 6'b010101;
12'b11101111100010: data = 6'b010101;
12'b11101111100011: data = 6'b010101;
12'b11101111100100: data = 6'b010101;
12'b11101111100101: data = 6'b010101;
12'b11101111100110: data = 6'b010101;
12'b11101111100111: data = 6'b010101;
12'b11101111101000: data = 6'b010101;
12'b11101111101001: data = 6'b010101;
12'b11101111101010: data = 6'b010101;
12'b11101111101011: data = 6'b010101;
12'b11101111101100: data = 6'b010101;
12'b11101111101101: data = 6'b010101;
12'b11101111101110: data = 6'b010101;
12'b11101111101111: data = 6'b010101;
12'b11101111110000: data = 6'b010101;
12'b11101111110001: data = 6'b010101;
12'b11101111110010: data = 6'b010101;
12'b11101111110011: data = 6'b010101;
12'b11101111110100: data = 6'b010101;
12'b11101111110101: data = 6'b010101;
12'b11101111110110: data = 6'b010101;
12'b11101111110111: data = 6'b010101;
12'b11101111111000: data = 6'b010101;
12'b11101111111001: data = 6'b000000;
12'b11101111111010: data = 6'b010101;
12'b11101111111011: data = 6'b000000;
12'b11101111111100: data = 6'b000000;
12'b11101111111101: data = 6'b000000;
12'b11101111111110: data = 6'b000000;
12'b11101111111111: data = 6'b000000;
12'b111011110000000: data = 6'b000000;
12'b111011110000001: data = 6'b000000;
12'b111011110000010: data = 6'b000000;
12'b111011110000011: data = 6'b000000;
12'b111011110000100: data = 6'b000000;
12'b111011110000101: data = 6'b000000;
12'b111011110000110: data = 6'b000000;
12'b111011110000111: data = 6'b000000;
12'b111011110001000: data = 6'b000000;
12'b111011110001001: data = 6'b000000;
12'b111011110001010: data = 6'b000000;
12'b111011110001011: data = 6'b000000;
12'b111011110001100: data = 6'b000000;
12'b111011110001101: data = 6'b000000;
12'b111011110001110: data = 6'b101010;
12'b111011110001111: data = 6'b101010;
12'b111011110010000: data = 6'b101010;
12'b111011110010001: data = 6'b101010;
12'b111011110010010: data = 6'b010101;
12'b111011110010011: data = 6'b010101;
12'b111011110010100: data = 6'b010101;
12'b111011110010101: data = 6'b010101;
12'b111011110010110: data = 6'b010101;
12'b111011110010111: data = 6'b010101;
12'b111011110011000: data = 6'b010101;
12'b111011110011001: data = 6'b010101;
12'b111011110011010: data = 6'b010101;
12'b111011110011011: data = 6'b010101;
12'b111011110011100: data = 6'b010101;
12'b111011110011101: data = 6'b010101;
12'b111011110011110: data = 6'b010101;
12'b111011110011111: data = 6'b010101;
12'b111011110100000: data = 6'b010101;
12'b111011110100001: data = 6'b010101;
12'b111011110100010: data = 6'b010101;
12'b111011110100011: data = 6'b010101;
12'b111011110100100: data = 6'b010101;
12'b111011110100101: data = 6'b010101;
12'b111011110100110: data = 6'b010101;
12'b111011110100111: data = 6'b010101;
12'b111011110101000: data = 6'b010101;
12'b111011110101001: data = 6'b010101;
12'b111011110101010: data = 6'b010101;
12'b1111000000000: data = 6'b010101;
12'b1111000000001: data = 6'b010101;
12'b1111000000010: data = 6'b010101;
12'b1111000000011: data = 6'b010101;
12'b1111000000100: data = 6'b010101;
12'b1111000000101: data = 6'b010101;
12'b1111000000110: data = 6'b010101;
12'b1111000000111: data = 6'b010101;
12'b1111000001000: data = 6'b010101;
12'b1111000001001: data = 6'b010101;
12'b1111000001010: data = 6'b010101;
12'b1111000001011: data = 6'b010101;
12'b1111000001100: data = 6'b010101;
12'b1111000001101: data = 6'b010101;
12'b1111000001110: data = 6'b010101;
12'b1111000001111: data = 6'b010101;
12'b1111000010000: data = 6'b010101;
12'b1111000010001: data = 6'b010101;
12'b1111000010010: data = 6'b010101;
12'b1111000010011: data = 6'b010101;
12'b1111000010100: data = 6'b010101;
12'b1111000010101: data = 6'b010101;
12'b1111000010110: data = 6'b010101;
12'b1111000010111: data = 6'b010101;
12'b1111000011000: data = 6'b010101;
12'b1111000011001: data = 6'b101010;
12'b1111000011010: data = 6'b101010;
12'b1111000011011: data = 6'b101010;
12'b1111000011100: data = 6'b101010;
12'b1111000011101: data = 6'b101010;
12'b1111000011110: data = 6'b101010;
12'b1111000011111: data = 6'b101010;
12'b1111000100000: data = 6'b101010;
12'b1111000100001: data = 6'b101010;
12'b1111000100010: data = 6'b010101;
12'b1111000100011: data = 6'b010101;
12'b1111000100100: data = 6'b010101;
12'b1111000100101: data = 6'b010101;
12'b1111000100110: data = 6'b010101;
12'b1111000100111: data = 6'b010101;
12'b1111000101000: data = 6'b010101;
12'b1111000101001: data = 6'b010101;
12'b1111000101010: data = 6'b010101;
12'b1111000101011: data = 6'b010101;
12'b1111000101100: data = 6'b010101;
12'b1111000101101: data = 6'b010101;
12'b1111000101110: data = 6'b010101;
12'b1111000101111: data = 6'b010101;
12'b1111000110000: data = 6'b010101;
12'b1111000110001: data = 6'b010101;
12'b1111000110010: data = 6'b010101;
12'b1111000110011: data = 6'b010101;
12'b1111000110100: data = 6'b010101;
12'b1111000110101: data = 6'b010101;
12'b1111000110110: data = 6'b010101;
12'b1111000110111: data = 6'b010101;
12'b1111000111000: data = 6'b010101;
12'b1111000111001: data = 6'b010101;
12'b1111000111010: data = 6'b010101;
12'b1111000111011: data = 6'b010101;
12'b1111000111100: data = 6'b010101;
12'b1111000111101: data = 6'b010101;
12'b1111000111110: data = 6'b010101;
12'b1111000111111: data = 6'b010101;
12'b11110001000000: data = 6'b010101;
12'b11110001000001: data = 6'b010101;
12'b11110001000010: data = 6'b010101;
12'b11110001000011: data = 6'b010101;
12'b11110001000100: data = 6'b010101;
12'b11110001000101: data = 6'b010101;
12'b11110001000110: data = 6'b010101;
12'b11110001000111: data = 6'b010101;
12'b11110001001000: data = 6'b010101;
12'b11110001001001: data = 6'b010101;
12'b11110001001010: data = 6'b010101;
12'b11110001001011: data = 6'b010101;
12'b11110001001100: data = 6'b010101;
12'b11110001001101: data = 6'b010101;
12'b11110001001110: data = 6'b010101;
12'b11110001001111: data = 6'b010101;
12'b11110001010000: data = 6'b010101;
12'b11110001010001: data = 6'b010101;
12'b11110001010010: data = 6'b010101;
12'b11110001010011: data = 6'b010101;
12'b11110001010100: data = 6'b010101;
12'b11110001010101: data = 6'b010101;
12'b11110001010110: data = 6'b010101;
12'b11110001010111: data = 6'b010101;
12'b11110001011000: data = 6'b010101;
12'b11110001011001: data = 6'b010101;
12'b11110001011010: data = 6'b010101;
12'b11110001011011: data = 6'b010101;
12'b11110001011100: data = 6'b010101;
12'b11110001011101: data = 6'b010101;
12'b11110001011110: data = 6'b010101;
12'b11110001011111: data = 6'b010101;
12'b11110001100000: data = 6'b010101;
12'b11110001100001: data = 6'b010101;
12'b11110001100010: data = 6'b010101;
12'b11110001100011: data = 6'b010101;
12'b11110001100100: data = 6'b010101;
12'b11110001100101: data = 6'b010101;
12'b11110001100110: data = 6'b010101;
12'b11110001100111: data = 6'b010101;
12'b11110001101000: data = 6'b010101;
12'b11110001101001: data = 6'b010101;
12'b11110001101010: data = 6'b010101;
12'b11110001101011: data = 6'b010101;
12'b11110001101100: data = 6'b010101;
12'b11110001101101: data = 6'b010101;
12'b11110001101110: data = 6'b010101;
12'b11110001101111: data = 6'b010101;
12'b11110001110000: data = 6'b010101;
12'b11110001110001: data = 6'b010101;
12'b11110001110010: data = 6'b010101;
12'b11110001110011: data = 6'b010101;
12'b11110001110100: data = 6'b010101;
12'b11110001110101: data = 6'b010101;
12'b11110001110110: data = 6'b010101;
12'b11110001110111: data = 6'b010101;
12'b11110001111000: data = 6'b010101;
12'b11110001111001: data = 6'b010101;
12'b11110001111010: data = 6'b010101;
12'b11110001111011: data = 6'b010101;
12'b11110001111100: data = 6'b010101;
12'b11110001111101: data = 6'b010101;
12'b11110001111110: data = 6'b010101;
12'b11110001111111: data = 6'b010101;
12'b111100010000000: data = 6'b010101;
12'b111100010000001: data = 6'b010101;
12'b111100010000010: data = 6'b010101;
12'b111100010000011: data = 6'b010101;
12'b111100010000100: data = 6'b010101;
12'b111100010000101: data = 6'b010101;
12'b111100010000110: data = 6'b010101;
12'b111100010000111: data = 6'b010101;
12'b111100010001000: data = 6'b010101;
12'b111100010001001: data = 6'b010101;
12'b111100010001010: data = 6'b010101;
12'b111100010001011: data = 6'b101010;
12'b111100010001100: data = 6'b101010;
12'b111100010001101: data = 6'b101010;
12'b111100010001110: data = 6'b101010;
12'b111100010001111: data = 6'b101010;
12'b111100010010000: data = 6'b101010;
12'b111100010010001: data = 6'b101010;
12'b111100010010010: data = 6'b010101;
12'b111100010010011: data = 6'b010101;
12'b111100010010100: data = 6'b010101;
12'b111100010010101: data = 6'b010101;
12'b111100010010110: data = 6'b010101;
12'b111100010010111: data = 6'b010101;
12'b111100010011000: data = 6'b010101;
12'b111100010011001: data = 6'b010101;
12'b111100010011010: data = 6'b010101;
12'b111100010011011: data = 6'b010101;
12'b111100010011100: data = 6'b010101;
12'b111100010011101: data = 6'b010101;
12'b111100010011110: data = 6'b010101;
12'b111100010011111: data = 6'b010101;
12'b111100010100000: data = 6'b010101;
12'b111100010100001: data = 6'b010101;
12'b111100010100010: data = 6'b010101;
12'b111100010100011: data = 6'b010101;
12'b111100010100100: data = 6'b010101;
12'b111100010100101: data = 6'b010101;
12'b111100010100110: data = 6'b010101;
12'b111100010100111: data = 6'b010101;
12'b111100010101000: data = 6'b010101;
12'b111100010101001: data = 6'b010101;
12'b111100010101010: data = 6'b010101;
12'b1111001000000: data = 6'b010101;
12'b1111001000001: data = 6'b010101;
12'b1111001000010: data = 6'b010101;
12'b1111001000011: data = 6'b010101;
12'b1111001000100: data = 6'b010101;
12'b1111001000101: data = 6'b010101;
12'b1111001000110: data = 6'b010101;
12'b1111001000111: data = 6'b010101;
12'b1111001001000: data = 6'b010101;
12'b1111001001001: data = 6'b010101;
12'b1111001001010: data = 6'b010101;
12'b1111001001011: data = 6'b010101;
12'b1111001001100: data = 6'b010101;
12'b1111001001101: data = 6'b010101;
12'b1111001001110: data = 6'b010101;
12'b1111001001111: data = 6'b010101;
12'b1111001010000: data = 6'b010101;
12'b1111001010001: data = 6'b010101;
12'b1111001010010: data = 6'b010101;
12'b1111001010011: data = 6'b010101;
12'b1111001010100: data = 6'b010101;
12'b1111001010101: data = 6'b010101;
12'b1111001010110: data = 6'b010101;
12'b1111001010111: data = 6'b010101;
12'b1111001011000: data = 6'b010101;
12'b1111001011001: data = 6'b101010;
12'b1111001011010: data = 6'b101010;
12'b1111001011011: data = 6'b101010;
12'b1111001011100: data = 6'b101010;
12'b1111001011101: data = 6'b101010;
12'b1111001011110: data = 6'b101010;
12'b1111001011111: data = 6'b101010;
12'b1111001100000: data = 6'b101010;
12'b1111001100001: data = 6'b101010;
12'b1111001100010: data = 6'b101010;
12'b1111001100011: data = 6'b010101;
12'b1111001100100: data = 6'b010101;
12'b1111001100101: data = 6'b010101;
12'b1111001100110: data = 6'b010101;
12'b1111001100111: data = 6'b010101;
12'b1111001101000: data = 6'b010101;
12'b1111001101001: data = 6'b010101;
12'b1111001101010: data = 6'b010101;
12'b1111001101011: data = 6'b010101;
12'b1111001101100: data = 6'b010101;
12'b1111001101101: data = 6'b010101;
12'b1111001101110: data = 6'b010101;
12'b1111001101111: data = 6'b010101;
12'b1111001110000: data = 6'b010101;
12'b1111001110001: data = 6'b010101;
12'b1111001110010: data = 6'b010101;
12'b1111001110011: data = 6'b010101;
12'b1111001110100: data = 6'b010101;
12'b1111001110101: data = 6'b010101;
12'b1111001110110: data = 6'b010101;
12'b1111001110111: data = 6'b010101;
12'b1111001111000: data = 6'b010101;
12'b1111001111001: data = 6'b010101;
12'b1111001111010: data = 6'b010101;
12'b1111001111011: data = 6'b010101;
12'b1111001111100: data = 6'b010101;
12'b1111001111101: data = 6'b010101;
12'b1111001111110: data = 6'b010101;
12'b1111001111111: data = 6'b010101;
12'b11110011000000: data = 6'b010101;
12'b11110011000001: data = 6'b010101;
12'b11110011000010: data = 6'b010101;
12'b11110011000011: data = 6'b010101;
12'b11110011000100: data = 6'b010101;
12'b11110011000101: data = 6'b010101;
12'b11110011000110: data = 6'b010101;
12'b11110011000111: data = 6'b010101;
12'b11110011001000: data = 6'b010101;
12'b11110011001001: data = 6'b010101;
12'b11110011001010: data = 6'b010101;
12'b11110011001011: data = 6'b010101;
12'b11110011001100: data = 6'b010101;
12'b11110011001101: data = 6'b010101;
12'b11110011001110: data = 6'b010101;
12'b11110011001111: data = 6'b010101;
12'b11110011010000: data = 6'b010101;
12'b11110011010001: data = 6'b010101;
12'b11110011010010: data = 6'b010101;
12'b11110011010011: data = 6'b010101;
12'b11110011010100: data = 6'b010101;
12'b11110011010101: data = 6'b010101;
12'b11110011010110: data = 6'b010101;
12'b11110011010111: data = 6'b010101;
12'b11110011011000: data = 6'b010101;
12'b11110011011001: data = 6'b010101;
12'b11110011011010: data = 6'b010101;
12'b11110011011011: data = 6'b010101;
12'b11110011011100: data = 6'b010101;
12'b11110011011101: data = 6'b010101;
12'b11110011011110: data = 6'b010101;
12'b11110011011111: data = 6'b010101;
12'b11110011100000: data = 6'b010101;
12'b11110011100001: data = 6'b010101;
12'b11110011100010: data = 6'b010101;
12'b11110011100011: data = 6'b010101;
12'b11110011100100: data = 6'b010101;
12'b11110011100101: data = 6'b010101;
12'b11110011100110: data = 6'b010101;
12'b11110011100111: data = 6'b010101;
12'b11110011101000: data = 6'b010101;
12'b11110011101001: data = 6'b010101;
12'b11110011101010: data = 6'b010101;
12'b11110011101011: data = 6'b010101;
12'b11110011101100: data = 6'b010101;
12'b11110011101101: data = 6'b010101;
12'b11110011101110: data = 6'b010101;
12'b11110011101111: data = 6'b010101;
12'b11110011110000: data = 6'b010101;
12'b11110011110001: data = 6'b010101;
12'b11110011110010: data = 6'b010101;
12'b11110011110011: data = 6'b010101;
12'b11110011110100: data = 6'b010101;
12'b11110011110101: data = 6'b010101;
12'b11110011110110: data = 6'b010101;
12'b11110011110111: data = 6'b010101;
12'b11110011111000: data = 6'b010101;
12'b11110011111001: data = 6'b010101;
12'b11110011111010: data = 6'b010101;
12'b11110011111011: data = 6'b010101;
12'b11110011111100: data = 6'b010101;
12'b11110011111101: data = 6'b010101;
12'b11110011111110: data = 6'b010101;
12'b11110011111111: data = 6'b010101;
12'b111100110000000: data = 6'b010101;
12'b111100110000001: data = 6'b010101;
12'b111100110000010: data = 6'b010101;
12'b111100110000011: data = 6'b010101;
12'b111100110000100: data = 6'b010101;
12'b111100110000101: data = 6'b010101;
12'b111100110000110: data = 6'b010101;
12'b111100110000111: data = 6'b010101;
12'b111100110001000: data = 6'b010101;
12'b111100110001001: data = 6'b101010;
12'b111100110001010: data = 6'b101010;
12'b111100110001011: data = 6'b101010;
12'b111100110001100: data = 6'b111110;
12'b111100110001101: data = 6'b101010;
12'b111100110001110: data = 6'b101010;
12'b111100110001111: data = 6'b101010;
12'b111100110010000: data = 6'b101010;
12'b111100110010001: data = 6'b101010;
12'b111100110010010: data = 6'b010101;
12'b111100110010011: data = 6'b010101;
12'b111100110010100: data = 6'b010101;
12'b111100110010101: data = 6'b010101;
12'b111100110010110: data = 6'b010101;
12'b111100110010111: data = 6'b010101;
12'b111100110011000: data = 6'b010101;
12'b111100110011001: data = 6'b010101;
12'b111100110011010: data = 6'b010101;
12'b111100110011011: data = 6'b010101;
12'b111100110011100: data = 6'b010101;
12'b111100110011101: data = 6'b010101;
12'b111100110011110: data = 6'b010101;
12'b111100110011111: data = 6'b010101;
12'b111100110100000: data = 6'b010101;
12'b111100110100001: data = 6'b010101;
12'b111100110100010: data = 6'b010101;
12'b111100110100011: data = 6'b010101;
12'b111100110100100: data = 6'b010101;
12'b111100110100101: data = 6'b010101;
12'b111100110100110: data = 6'b010101;
12'b111100110100111: data = 6'b010101;
12'b111100110101000: data = 6'b010101;
12'b111100110101001: data = 6'b010101;
12'b111100110101010: data = 6'b010101;
12'b1111010000000: data = 6'b010101;
12'b1111010000001: data = 6'b010101;
12'b1111010000010: data = 6'b010101;
12'b1111010000011: data = 6'b010101;
12'b1111010000100: data = 6'b010101;
12'b1111010000101: data = 6'b010101;
12'b1111010000110: data = 6'b010101;
12'b1111010000111: data = 6'b010101;
12'b1111010001000: data = 6'b010101;
12'b1111010001001: data = 6'b010101;
12'b1111010001010: data = 6'b010101;
12'b1111010001011: data = 6'b010101;
12'b1111010001100: data = 6'b010101;
12'b1111010001101: data = 6'b010101;
12'b1111010001110: data = 6'b010101;
12'b1111010001111: data = 6'b010101;
12'b1111010010000: data = 6'b010101;
12'b1111010010001: data = 6'b010101;
12'b1111010010010: data = 6'b010101;
12'b1111010010011: data = 6'b010101;
12'b1111010010100: data = 6'b010101;
12'b1111010010101: data = 6'b010101;
12'b1111010010110: data = 6'b010101;
12'b1111010010111: data = 6'b010101;
12'b1111010011000: data = 6'b010101;
12'b1111010011001: data = 6'b010101;
12'b1111010011010: data = 6'b101010;
12'b1111010011011: data = 6'b101010;
12'b1111010011100: data = 6'b101010;
12'b1111010011101: data = 6'b101010;
12'b1111010011110: data = 6'b101010;
12'b1111010011111: data = 6'b101010;
12'b1111010100000: data = 6'b101010;
12'b1111010100001: data = 6'b101010;
12'b1111010100010: data = 6'b101010;
12'b1111010100011: data = 6'b101001;
12'b1111010100100: data = 6'b010101;
12'b1111010100101: data = 6'b010101;
12'b1111010100110: data = 6'b010101;
12'b1111010100111: data = 6'b010101;
12'b1111010101000: data = 6'b010101;
12'b1111010101001: data = 6'b010101;
12'b1111010101010: data = 6'b010101;
12'b1111010101011: data = 6'b010101;
12'b1111010101100: data = 6'b010101;
12'b1111010101101: data = 6'b010101;
12'b1111010101110: data = 6'b010101;
12'b1111010101111: data = 6'b010101;
12'b1111010110000: data = 6'b010101;
12'b1111010110001: data = 6'b010101;
12'b1111010110010: data = 6'b010101;
12'b1111010110011: data = 6'b010101;
12'b1111010110100: data = 6'b010101;
12'b1111010110101: data = 6'b010101;
12'b1111010110110: data = 6'b010101;
12'b1111010110111: data = 6'b010101;
12'b1111010111000: data = 6'b010101;
12'b1111010111001: data = 6'b010101;
12'b1111010111010: data = 6'b010101;
12'b1111010111011: data = 6'b010101;
12'b1111010111100: data = 6'b010101;
12'b1111010111101: data = 6'b010101;
12'b1111010111110: data = 6'b010101;
12'b1111010111111: data = 6'b010101;
12'b11110101000000: data = 6'b010101;
12'b11110101000001: data = 6'b010101;
12'b11110101000010: data = 6'b010101;
12'b11110101000011: data = 6'b010101;
12'b11110101000100: data = 6'b010101;
12'b11110101000101: data = 6'b010101;
12'b11110101000110: data = 6'b010101;
12'b11110101000111: data = 6'b010101;
12'b11110101001000: data = 6'b010101;
12'b11110101001001: data = 6'b010101;
12'b11110101001010: data = 6'b010101;
12'b11110101001011: data = 6'b010101;
12'b11110101001100: data = 6'b010101;
12'b11110101001101: data = 6'b010101;
12'b11110101001110: data = 6'b010101;
12'b11110101001111: data = 6'b010101;
12'b11110101010000: data = 6'b010101;
12'b11110101010001: data = 6'b010101;
12'b11110101010010: data = 6'b010101;
12'b11110101010011: data = 6'b010101;
12'b11110101010100: data = 6'b010101;
12'b11110101010101: data = 6'b010101;
12'b11110101010110: data = 6'b010101;
12'b11110101010111: data = 6'b010101;
12'b11110101011000: data = 6'b010101;
12'b11110101011001: data = 6'b010101;
12'b11110101011010: data = 6'b010101;
12'b11110101011011: data = 6'b010101;
12'b11110101011100: data = 6'b010101;
12'b11110101011101: data = 6'b010101;
12'b11110101011110: data = 6'b010101;
12'b11110101011111: data = 6'b010101;
12'b11110101100000: data = 6'b010101;
12'b11110101100001: data = 6'b010101;
12'b11110101100010: data = 6'b010101;
12'b11110101100011: data = 6'b010101;
12'b11110101100100: data = 6'b010101;
12'b11110101100101: data = 6'b010101;
12'b11110101100110: data = 6'b010101;
12'b11110101100111: data = 6'b010101;
12'b11110101101000: data = 6'b010101;
12'b11110101101001: data = 6'b010101;
12'b11110101101010: data = 6'b010101;
12'b11110101101011: data = 6'b010101;
12'b11110101101100: data = 6'b010101;
12'b11110101101101: data = 6'b010101;
12'b11110101101110: data = 6'b010101;
12'b11110101101111: data = 6'b010101;
12'b11110101110000: data = 6'b010101;
12'b11110101110001: data = 6'b010101;
12'b11110101110010: data = 6'b010101;
12'b11110101110011: data = 6'b010101;
12'b11110101110100: data = 6'b010101;
12'b11110101110101: data = 6'b010101;
12'b11110101110110: data = 6'b010101;
12'b11110101110111: data = 6'b010101;
12'b11110101111000: data = 6'b010101;
12'b11110101111001: data = 6'b010101;
12'b11110101111010: data = 6'b010101;
12'b11110101111011: data = 6'b010101;
12'b11110101111100: data = 6'b010101;
12'b11110101111101: data = 6'b010101;
12'b11110101111110: data = 6'b010101;
12'b11110101111111: data = 6'b010101;
12'b111101010000000: data = 6'b010101;
12'b111101010000001: data = 6'b010101;
12'b111101010000010: data = 6'b010101;
12'b111101010000011: data = 6'b010101;
12'b111101010000100: data = 6'b010101;
12'b111101010000101: data = 6'b010101;
12'b111101010000110: data = 6'b010101;
12'b111101010000111: data = 6'b100101;
12'b111101010001000: data = 6'b101010;
12'b111101010001001: data = 6'b101010;
12'b111101010001010: data = 6'b101010;
12'b111101010001011: data = 6'b101010;
12'b111101010001100: data = 6'b101010;
12'b111101010001101: data = 6'b101010;
12'b111101010001110: data = 6'b101010;
12'b111101010001111: data = 6'b101010;
12'b111101010010000: data = 6'b101010;
12'b111101010010001: data = 6'b010101;
12'b111101010010010: data = 6'b010101;
12'b111101010010011: data = 6'b010101;
12'b111101010010100: data = 6'b010101;
12'b111101010010101: data = 6'b010101;
12'b111101010010110: data = 6'b010101;
12'b111101010010111: data = 6'b010101;
12'b111101010011000: data = 6'b010101;
12'b111101010011001: data = 6'b010101;
12'b111101010011010: data = 6'b010101;
12'b111101010011011: data = 6'b010101;
12'b111101010011100: data = 6'b010101;
12'b111101010011101: data = 6'b010101;
12'b111101010011110: data = 6'b010101;
12'b111101010011111: data = 6'b010101;
12'b111101010100000: data = 6'b010101;
12'b111101010100001: data = 6'b010101;
12'b111101010100010: data = 6'b010101;
12'b111101010100011: data = 6'b010101;
12'b111101010100100: data = 6'b010101;
12'b111101010100101: data = 6'b010101;
12'b111101010100110: data = 6'b010101;
12'b111101010100111: data = 6'b010101;
12'b111101010101000: data = 6'b010101;
12'b111101010101001: data = 6'b010101;
12'b111101010101010: data = 6'b010101;
12'b1111011000000: data = 6'b010101;
12'b1111011000001: data = 6'b010101;
12'b1111011000010: data = 6'b010101;
12'b1111011000011: data = 6'b010101;
12'b1111011000100: data = 6'b010101;
12'b1111011000101: data = 6'b010101;
12'b1111011000110: data = 6'b010101;
12'b1111011000111: data = 6'b010101;
12'b1111011001000: data = 6'b010101;
12'b1111011001001: data = 6'b010101;
12'b1111011001010: data = 6'b010101;
12'b1111011001011: data = 6'b010101;
12'b1111011001100: data = 6'b010101;
12'b1111011001101: data = 6'b010101;
12'b1111011001110: data = 6'b010101;
12'b1111011001111: data = 6'b010101;
12'b1111011010000: data = 6'b010101;
12'b1111011010001: data = 6'b010101;
12'b1111011010010: data = 6'b010101;
12'b1111011010011: data = 6'b010101;
12'b1111011010100: data = 6'b010101;
12'b1111011010101: data = 6'b010101;
12'b1111011010110: data = 6'b010101;
12'b1111011010111: data = 6'b010101;
12'b1111011011000: data = 6'b010101;
12'b1111011011001: data = 6'b010101;
12'b1111011011010: data = 6'b101010;
12'b1111011011011: data = 6'b101010;
12'b1111011011100: data = 6'b101010;
12'b1111011011101: data = 6'b101010;
12'b1111011011110: data = 6'b101010;
12'b1111011011111: data = 6'b101010;
12'b1111011100000: data = 6'b101010;
12'b1111011100001: data = 6'b101010;
12'b1111011100010: data = 6'b101010;
12'b1111011100011: data = 6'b101010;
12'b1111011100100: data = 6'b101010;
12'b1111011100101: data = 6'b010101;
12'b1111011100110: data = 6'b010101;
12'b1111011100111: data = 6'b010101;
12'b1111011101000: data = 6'b010101;
12'b1111011101001: data = 6'b010101;
12'b1111011101010: data = 6'b010101;
12'b1111011101011: data = 6'b010101;
12'b1111011101100: data = 6'b010101;
12'b1111011101101: data = 6'b010101;
12'b1111011101110: data = 6'b010101;
12'b1111011101111: data = 6'b010101;
12'b1111011110000: data = 6'b010101;
12'b1111011110001: data = 6'b010101;
12'b1111011110010: data = 6'b010101;
12'b1111011110011: data = 6'b010101;
12'b1111011110100: data = 6'b010101;
12'b1111011110101: data = 6'b010101;
12'b1111011110110: data = 6'b010101;
12'b1111011110111: data = 6'b010101;
12'b1111011111000: data = 6'b010101;
12'b1111011111001: data = 6'b010101;
12'b1111011111010: data = 6'b010101;
12'b1111011111011: data = 6'b010101;
12'b1111011111100: data = 6'b010101;
12'b1111011111101: data = 6'b010101;
12'b1111011111110: data = 6'b010101;
12'b1111011111111: data = 6'b010101;
12'b11110111000000: data = 6'b010101;
12'b11110111000001: data = 6'b010101;
12'b11110111000010: data = 6'b010101;
12'b11110111000011: data = 6'b010101;
12'b11110111000100: data = 6'b010101;
12'b11110111000101: data = 6'b010101;
12'b11110111000110: data = 6'b010101;
12'b11110111000111: data = 6'b010101;
12'b11110111001000: data = 6'b010101;
12'b11110111001001: data = 6'b010101;
12'b11110111001010: data = 6'b010101;
12'b11110111001011: data = 6'b010101;
12'b11110111001100: data = 6'b010101;
12'b11110111001101: data = 6'b010101;
12'b11110111001110: data = 6'b010101;
12'b11110111001111: data = 6'b010101;
12'b11110111010000: data = 6'b010101;
12'b11110111010001: data = 6'b010101;
12'b11110111010010: data = 6'b010101;
12'b11110111010011: data = 6'b010101;
12'b11110111010100: data = 6'b010101;
12'b11110111010101: data = 6'b010101;
12'b11110111010110: data = 6'b010101;
12'b11110111010111: data = 6'b010101;
12'b11110111011000: data = 6'b010101;
12'b11110111011001: data = 6'b010101;
12'b11110111011010: data = 6'b010101;
12'b11110111011011: data = 6'b010101;
12'b11110111011100: data = 6'b010101;
12'b11110111011101: data = 6'b010101;
12'b11110111011110: data = 6'b010101;
12'b11110111011111: data = 6'b010101;
12'b11110111100000: data = 6'b010101;
12'b11110111100001: data = 6'b010101;
12'b11110111100010: data = 6'b010101;
12'b11110111100011: data = 6'b010101;
12'b11110111100100: data = 6'b010101;
12'b11110111100101: data = 6'b010101;
12'b11110111100110: data = 6'b010101;
12'b11110111100111: data = 6'b010101;
12'b11110111101000: data = 6'b010101;
12'b11110111101001: data = 6'b010101;
12'b11110111101010: data = 6'b010101;
12'b11110111101011: data = 6'b010101;
12'b11110111101100: data = 6'b010101;
12'b11110111101101: data = 6'b010101;
12'b11110111101110: data = 6'b010101;
12'b11110111101111: data = 6'b010101;
12'b11110111110000: data = 6'b010101;
12'b11110111110001: data = 6'b010101;
12'b11110111110010: data = 6'b010101;
12'b11110111110011: data = 6'b010101;
12'b11110111110100: data = 6'b010101;
12'b11110111110101: data = 6'b010101;
12'b11110111110110: data = 6'b010101;
12'b11110111110111: data = 6'b010101;
12'b11110111111000: data = 6'b010101;
12'b11110111111001: data = 6'b010101;
12'b11110111111010: data = 6'b010101;
12'b11110111111011: data = 6'b010101;
12'b11110111111100: data = 6'b010101;
12'b11110111111101: data = 6'b010101;
12'b11110111111110: data = 6'b010101;
12'b11110111111111: data = 6'b010101;
12'b111101110000000: data = 6'b010101;
12'b111101110000001: data = 6'b010101;
12'b111101110000010: data = 6'b010101;
12'b111101110000011: data = 6'b010101;
12'b111101110000100: data = 6'b010101;
12'b111101110000101: data = 6'b010101;
12'b111101110000110: data = 6'b100101;
12'b111101110000111: data = 6'b101010;
12'b111101110001000: data = 6'b101010;
12'b111101110001001: data = 6'b101010;
12'b111101110001010: data = 6'b101010;
12'b111101110001011: data = 6'b101010;
12'b111101110001100: data = 6'b101010;
12'b111101110001101: data = 6'b101010;
12'b111101110001110: data = 6'b101010;
12'b111101110001111: data = 6'b101010;
12'b111101110010000: data = 6'b101010;
12'b111101110010001: data = 6'b010101;
12'b111101110010010: data = 6'b010101;
12'b111101110010011: data = 6'b010101;
12'b111101110010100: data = 6'b010101;
12'b111101110010101: data = 6'b010101;
12'b111101110010110: data = 6'b010101;
12'b111101110010111: data = 6'b010101;
12'b111101110011000: data = 6'b010101;
12'b111101110011001: data = 6'b010101;
12'b111101110011010: data = 6'b010101;
12'b111101110011011: data = 6'b010101;
12'b111101110011100: data = 6'b010101;
12'b111101110011101: data = 6'b010101;
12'b111101110011110: data = 6'b010101;
12'b111101110011111: data = 6'b010101;
12'b111101110100000: data = 6'b010101;
12'b111101110100001: data = 6'b010101;
12'b111101110100010: data = 6'b010101;
12'b111101110100011: data = 6'b010101;
12'b111101110100100: data = 6'b010101;
12'b111101110100101: data = 6'b010101;
12'b111101110100110: data = 6'b010101;
12'b111101110100111: data = 6'b010101;
12'b111101110101000: data = 6'b010101;
12'b111101110101001: data = 6'b010101;
12'b111101110101010: data = 6'b010101;
12'b1111100000000: data = 6'b010101;
12'b1111100000001: data = 6'b010101;
12'b1111100000010: data = 6'b010101;
12'b1111100000011: data = 6'b010101;
12'b1111100000100: data = 6'b010101;
12'b1111100000101: data = 6'b010101;
12'b1111100000110: data = 6'b010101;
12'b1111100000111: data = 6'b010101;
12'b1111100001000: data = 6'b010101;
12'b1111100001001: data = 6'b010101;
12'b1111100001010: data = 6'b010101;
12'b1111100001011: data = 6'b010101;
12'b1111100001100: data = 6'b010101;
12'b1111100001101: data = 6'b010101;
12'b1111100001110: data = 6'b010101;
12'b1111100001111: data = 6'b010101;
12'b1111100010000: data = 6'b010101;
12'b1111100010001: data = 6'b010101;
12'b1111100010010: data = 6'b010101;
12'b1111100010011: data = 6'b010101;
12'b1111100010100: data = 6'b010101;
12'b1111100010101: data = 6'b010101;
12'b1111100010110: data = 6'b010101;
12'b1111100010111: data = 6'b010101;
12'b1111100011000: data = 6'b010101;
12'b1111100011001: data = 6'b010101;
12'b1111100011010: data = 6'b101010;
12'b1111100011011: data = 6'b101010;
12'b1111100011100: data = 6'b101010;
12'b1111100011101: data = 6'b101010;
12'b1111100011110: data = 6'b101010;
12'b1111100011111: data = 6'b101010;
12'b1111100100000: data = 6'b101010;
12'b1111100100001: data = 6'b101010;
12'b1111100100010: data = 6'b101010;
12'b1111100100011: data = 6'b101010;
12'b1111100100100: data = 6'b101010;
12'b1111100100101: data = 6'b010101;
12'b1111100100110: data = 6'b010101;
12'b1111100100111: data = 6'b010101;
12'b1111100101000: data = 6'b010101;
12'b1111100101001: data = 6'b010101;
12'b1111100101010: data = 6'b010101;
12'b1111100101011: data = 6'b010101;
12'b1111100101100: data = 6'b010101;
12'b1111100101101: data = 6'b010101;
12'b1111100101110: data = 6'b010101;
12'b1111100101111: data = 6'b010101;
12'b1111100110000: data = 6'b010101;
12'b1111100110001: data = 6'b010101;
12'b1111100110010: data = 6'b010101;
12'b1111100110011: data = 6'b010101;
12'b1111100110100: data = 6'b010101;
12'b1111100110101: data = 6'b010101;
12'b1111100110110: data = 6'b010101;
12'b1111100110111: data = 6'b010101;
12'b1111100111000: data = 6'b010101;
12'b1111100111001: data = 6'b010101;
12'b1111100111010: data = 6'b010101;
12'b1111100111011: data = 6'b010101;
12'b1111100111100: data = 6'b010101;
12'b1111100111101: data = 6'b010101;
12'b1111100111110: data = 6'b010101;
12'b1111100111111: data = 6'b010101;
12'b11111001000000: data = 6'b010101;
12'b11111001000001: data = 6'b010101;
12'b11111001000010: data = 6'b010101;
12'b11111001000011: data = 6'b010101;
12'b11111001000100: data = 6'b010101;
12'b11111001000101: data = 6'b010101;
12'b11111001000110: data = 6'b010101;
12'b11111001000111: data = 6'b010101;
12'b11111001001000: data = 6'b010101;
12'b11111001001001: data = 6'b010101;
12'b11111001001010: data = 6'b010101;
12'b11111001001011: data = 6'b010101;
12'b11111001001100: data = 6'b010101;
12'b11111001001101: data = 6'b010101;
12'b11111001001110: data = 6'b010101;
12'b11111001001111: data = 6'b010101;
12'b11111001010000: data = 6'b010101;
12'b11111001010001: data = 6'b010101;
12'b11111001010010: data = 6'b010101;
12'b11111001010011: data = 6'b010101;
12'b11111001010100: data = 6'b010101;
12'b11111001010101: data = 6'b010101;
12'b11111001010110: data = 6'b010101;
12'b11111001010111: data = 6'b010101;
12'b11111001011000: data = 6'b010101;
12'b11111001011001: data = 6'b010101;
12'b11111001011010: data = 6'b010101;
12'b11111001011011: data = 6'b010101;
12'b11111001011100: data = 6'b010101;
12'b11111001011101: data = 6'b010101;
12'b11111001011110: data = 6'b010101;
12'b11111001011111: data = 6'b010101;
12'b11111001100000: data = 6'b010101;
12'b11111001100001: data = 6'b010101;
12'b11111001100010: data = 6'b010101;
12'b11111001100011: data = 6'b010101;
12'b11111001100100: data = 6'b010101;
12'b11111001100101: data = 6'b010101;
12'b11111001100110: data = 6'b010101;
12'b11111001100111: data = 6'b010101;
12'b11111001101000: data = 6'b010101;
12'b11111001101001: data = 6'b010101;
12'b11111001101010: data = 6'b010101;
12'b11111001101011: data = 6'b010101;
12'b11111001101100: data = 6'b010101;
12'b11111001101101: data = 6'b010101;
12'b11111001101110: data = 6'b010101;
12'b11111001101111: data = 6'b010101;
12'b11111001110000: data = 6'b010101;
12'b11111001110001: data = 6'b010101;
12'b11111001110010: data = 6'b010101;
12'b11111001110011: data = 6'b010101;
12'b11111001110100: data = 6'b010101;
12'b11111001110101: data = 6'b010101;
12'b11111001110110: data = 6'b010101;
12'b11111001110111: data = 6'b010101;
12'b11111001111000: data = 6'b010101;
12'b11111001111001: data = 6'b010101;
12'b11111001111010: data = 6'b010101;
12'b11111001111011: data = 6'b010101;
12'b11111001111100: data = 6'b010101;
12'b11111001111101: data = 6'b010101;
12'b11111001111110: data = 6'b010101;
12'b11111001111111: data = 6'b010101;
12'b111110010000000: data = 6'b010101;
12'b111110010000001: data = 6'b010101;
12'b111110010000010: data = 6'b010101;
12'b111110010000011: data = 6'b010101;
12'b111110010000100: data = 6'b010101;
12'b111110010000101: data = 6'b010101;
12'b111110010000110: data = 6'b100101;
12'b111110010000111: data = 6'b101010;
12'b111110010001000: data = 6'b101010;
12'b111110010001001: data = 6'b101010;
12'b111110010001010: data = 6'b101010;
12'b111110010001011: data = 6'b101010;
12'b111110010001100: data = 6'b111010;
12'b111110010001101: data = 6'b101010;
12'b111110010001110: data = 6'b101010;
12'b111110010001111: data = 6'b101010;
12'b111110010010000: data = 6'b101010;
12'b111110010010001: data = 6'b010101;
12'b111110010010010: data = 6'b010101;
12'b111110010010011: data = 6'b010101;
12'b111110010010100: data = 6'b010101;
12'b111110010010101: data = 6'b010101;
12'b111110010010110: data = 6'b010101;
12'b111110010010111: data = 6'b010101;
12'b111110010011000: data = 6'b010101;
12'b111110010011001: data = 6'b010101;
12'b111110010011010: data = 6'b010101;
12'b111110010011011: data = 6'b010101;
12'b111110010011100: data = 6'b010101;
12'b111110010011101: data = 6'b010101;
12'b111110010011110: data = 6'b010101;
12'b111110010011111: data = 6'b010101;
12'b111110010100000: data = 6'b010101;
12'b111110010100001: data = 6'b010101;
12'b111110010100010: data = 6'b010101;
12'b111110010100011: data = 6'b010101;
12'b111110010100100: data = 6'b010101;
12'b111110010100101: data = 6'b010101;
12'b111110010100110: data = 6'b010101;
12'b111110010100111: data = 6'b010101;
12'b111110010101000: data = 6'b010101;
12'b111110010101001: data = 6'b010101;
12'b111110010101010: data = 6'b010101;
12'b1111101000000: data = 6'b010101;
12'b1111101000001: data = 6'b010101;
12'b1111101000010: data = 6'b010101;
12'b1111101000011: data = 6'b010101;
12'b1111101000100: data = 6'b010101;
12'b1111101000101: data = 6'b010101;
12'b1111101000110: data = 6'b010101;
12'b1111101000111: data = 6'b010101;
12'b1111101001000: data = 6'b010101;
12'b1111101001001: data = 6'b010101;
12'b1111101001010: data = 6'b010101;
12'b1111101001011: data = 6'b010101;
12'b1111101001100: data = 6'b010101;
12'b1111101001101: data = 6'b010101;
12'b1111101001110: data = 6'b010101;
12'b1111101001111: data = 6'b010101;
12'b1111101010000: data = 6'b010101;
12'b1111101010001: data = 6'b010101;
12'b1111101010010: data = 6'b010101;
12'b1111101010011: data = 6'b010101;
12'b1111101010100: data = 6'b010101;
12'b1111101010101: data = 6'b010101;
12'b1111101010110: data = 6'b010101;
12'b1111101010111: data = 6'b010101;
12'b1111101011000: data = 6'b010101;
12'b1111101011001: data = 6'b010101;
12'b1111101011010: data = 6'b101010;
12'b1111101011011: data = 6'b101010;
12'b1111101011100: data = 6'b101010;
12'b1111101011101: data = 6'b101010;
12'b1111101011110: data = 6'b101010;
12'b1111101011111: data = 6'b101010;
12'b1111101100000: data = 6'b101010;
12'b1111101100001: data = 6'b101010;
12'b1111101100010: data = 6'b101010;
12'b1111101100011: data = 6'b101010;
12'b1111101100100: data = 6'b101001;
12'b1111101100101: data = 6'b010101;
12'b1111101100110: data = 6'b010101;
12'b1111101100111: data = 6'b010101;
12'b1111101101000: data = 6'b010101;
12'b1111101101001: data = 6'b010101;
12'b1111101101010: data = 6'b010101;
12'b1111101101011: data = 6'b010101;
12'b1111101101100: data = 6'b010101;
12'b1111101101101: data = 6'b010101;
12'b1111101101110: data = 6'b010101;
12'b1111101101111: data = 6'b010101;
12'b1111101110000: data = 6'b010101;
12'b1111101110001: data = 6'b010101;
12'b1111101110010: data = 6'b010101;
12'b1111101110011: data = 6'b010101;
12'b1111101110100: data = 6'b010101;
12'b1111101110101: data = 6'b010101;
12'b1111101110110: data = 6'b010101;
12'b1111101110111: data = 6'b010101;
12'b1111101111000: data = 6'b010101;
12'b1111101111001: data = 6'b010101;
12'b1111101111010: data = 6'b010101;
12'b1111101111011: data = 6'b010101;
12'b1111101111100: data = 6'b010101;
12'b1111101111101: data = 6'b010101;
12'b1111101111110: data = 6'b010101;
12'b1111101111111: data = 6'b010101;
12'b11111011000000: data = 6'b010101;
12'b11111011000001: data = 6'b010101;
12'b11111011000010: data = 6'b010101;
12'b11111011000011: data = 6'b010101;
12'b11111011000100: data = 6'b010101;
12'b11111011000101: data = 6'b010101;
12'b11111011000110: data = 6'b010101;
12'b11111011000111: data = 6'b010101;
12'b11111011001000: data = 6'b010101;
12'b11111011001001: data = 6'b010101;
12'b11111011001010: data = 6'b010101;
12'b11111011001011: data = 6'b010101;
12'b11111011001100: data = 6'b010101;
12'b11111011001101: data = 6'b010101;
12'b11111011001110: data = 6'b010101;
12'b11111011001111: data = 6'b010101;
12'b11111011010000: data = 6'b010101;
12'b11111011010001: data = 6'b010101;
12'b11111011010010: data = 6'b010101;
12'b11111011010011: data = 6'b010101;
12'b11111011010100: data = 6'b010101;
12'b11111011010101: data = 6'b010101;
12'b11111011010110: data = 6'b010101;
12'b11111011010111: data = 6'b010101;
12'b11111011011000: data = 6'b010101;
12'b11111011011001: data = 6'b010101;
12'b11111011011010: data = 6'b010101;
12'b11111011011011: data = 6'b010101;
12'b11111011011100: data = 6'b010101;
12'b11111011011101: data = 6'b010101;
12'b11111011011110: data = 6'b010101;
12'b11111011011111: data = 6'b010101;
12'b11111011100000: data = 6'b010101;
12'b11111011100001: data = 6'b010101;
12'b11111011100010: data = 6'b010101;
12'b11111011100011: data = 6'b010101;
12'b11111011100100: data = 6'b010101;
12'b11111011100101: data = 6'b010101;
12'b11111011100110: data = 6'b010101;
12'b11111011100111: data = 6'b010101;
12'b11111011101000: data = 6'b010101;
12'b11111011101001: data = 6'b010101;
12'b11111011101010: data = 6'b010101;
12'b11111011101011: data = 6'b010101;
12'b11111011101100: data = 6'b010101;
12'b11111011101101: data = 6'b010101;
12'b11111011101110: data = 6'b010101;
12'b11111011101111: data = 6'b010101;
12'b11111011110000: data = 6'b010101;
12'b11111011110001: data = 6'b010101;
12'b11111011110010: data = 6'b010101;
12'b11111011110011: data = 6'b010101;
12'b11111011110100: data = 6'b010101;
12'b11111011110101: data = 6'b010101;
12'b11111011110110: data = 6'b010101;
12'b11111011110111: data = 6'b010101;
12'b11111011111000: data = 6'b010101;
12'b11111011111001: data = 6'b010101;
12'b11111011111010: data = 6'b010101;
12'b11111011111011: data = 6'b010101;
12'b11111011111100: data = 6'b010101;
12'b11111011111101: data = 6'b010101;
12'b11111011111110: data = 6'b010101;
12'b11111011111111: data = 6'b010101;
12'b111110110000000: data = 6'b010101;
12'b111110110000001: data = 6'b010101;
12'b111110110000010: data = 6'b010101;
12'b111110110000011: data = 6'b010101;
12'b111110110000100: data = 6'b010101;
12'b111110110000101: data = 6'b010101;
12'b111110110000110: data = 6'b101001;
12'b111110110000111: data = 6'b101001;
12'b111110110001000: data = 6'b101010;
12'b111110110001001: data = 6'b101010;
12'b111110110001010: data = 6'b101010;
12'b111110110001011: data = 6'b101010;
12'b111110110001100: data = 6'b101010;
12'b111110110001101: data = 6'b101010;
12'b111110110001110: data = 6'b101010;
12'b111110110001111: data = 6'b101010;
12'b111110110010000: data = 6'b101010;
12'b111110110010001: data = 6'b010101;
12'b111110110010010: data = 6'b010101;
12'b111110110010011: data = 6'b010101;
12'b111110110010100: data = 6'b010101;
12'b111110110010101: data = 6'b010101;
12'b111110110010110: data = 6'b010101;
12'b111110110010111: data = 6'b010101;
12'b111110110011000: data = 6'b010101;
12'b111110110011001: data = 6'b010101;
12'b111110110011010: data = 6'b010101;
12'b111110110011011: data = 6'b010101;
12'b111110110011100: data = 6'b010101;
12'b111110110011101: data = 6'b010101;
12'b111110110011110: data = 6'b010101;
12'b111110110011111: data = 6'b010101;
12'b111110110100000: data = 6'b010101;
12'b111110110100001: data = 6'b010101;
12'b111110110100010: data = 6'b010101;
12'b111110110100011: data = 6'b010101;
12'b111110110100100: data = 6'b010101;
12'b111110110100101: data = 6'b010101;
12'b111110110100110: data = 6'b010101;
12'b111110110100111: data = 6'b010101;
12'b111110110101000: data = 6'b010101;
12'b111110110101001: data = 6'b010101;
12'b111110110101010: data = 6'b010101;
12'b1111110000000: data = 6'b010101;
12'b1111110000001: data = 6'b010101;
12'b1111110000010: data = 6'b010101;
12'b1111110000011: data = 6'b010101;
12'b1111110000100: data = 6'b010101;
12'b1111110000101: data = 6'b010101;
12'b1111110000110: data = 6'b010101;
12'b1111110000111: data = 6'b010101;
12'b1111110001000: data = 6'b010101;
12'b1111110001001: data = 6'b010101;
12'b1111110001010: data = 6'b010101;
12'b1111110001011: data = 6'b010101;
12'b1111110001100: data = 6'b010101;
12'b1111110001101: data = 6'b010101;
12'b1111110001110: data = 6'b010101;
12'b1111110001111: data = 6'b010101;
12'b1111110010000: data = 6'b010101;
12'b1111110010001: data = 6'b010101;
12'b1111110010010: data = 6'b010101;
12'b1111110010011: data = 6'b010101;
12'b1111110010100: data = 6'b010101;
12'b1111110010101: data = 6'b010101;
12'b1111110010110: data = 6'b010101;
12'b1111110010111: data = 6'b010101;
12'b1111110011000: data = 6'b010101;
12'b1111110011001: data = 6'b010101;
12'b1111110011010: data = 6'b101010;
12'b1111110011011: data = 6'b101010;
12'b1111110011100: data = 6'b101010;
12'b1111110011101: data = 6'b010101;
12'b1111110011110: data = 6'b010101;
12'b1111110011111: data = 6'b010101;
12'b1111110100000: data = 6'b010101;
12'b1111110100001: data = 6'b010101;
12'b1111110100010: data = 6'b010101;
12'b1111110100011: data = 6'b010101;
12'b1111110100100: data = 6'b010101;
12'b1111110100101: data = 6'b010101;
12'b1111110100110: data = 6'b010101;
12'b1111110100111: data = 6'b010101;
12'b1111110101000: data = 6'b010101;
12'b1111110101001: data = 6'b010101;
12'b1111110101010: data = 6'b000000;
12'b1111110101011: data = 6'b000000;
12'b1111110101100: data = 6'b010101;
12'b1111110101101: data = 6'b010101;
12'b1111110101110: data = 6'b010101;
12'b1111110101111: data = 6'b010101;
12'b1111110110000: data = 6'b010101;
12'b1111110110001: data = 6'b010101;
12'b1111110110010: data = 6'b010101;
12'b1111110110011: data = 6'b010101;
12'b1111110110100: data = 6'b010101;
12'b1111110110101: data = 6'b010101;
12'b1111110110110: data = 6'b010101;
12'b1111110110111: data = 6'b010101;
12'b1111110111000: data = 6'b010101;
12'b1111110111001: data = 6'b010101;
12'b1111110111010: data = 6'b010101;
12'b1111110111011: data = 6'b010101;
12'b1111110111100: data = 6'b101010;
12'b1111110111101: data = 6'b101010;
12'b1111110111110: data = 6'b101010;
12'b1111110111111: data = 6'b010101;
12'b11111101000000: data = 6'b010101;
12'b11111101000001: data = 6'b010101;
12'b11111101000010: data = 6'b010101;
12'b11111101000011: data = 6'b010101;
12'b11111101000100: data = 6'b010101;
12'b11111101000101: data = 6'b010101;
12'b11111101000110: data = 6'b010101;
12'b11111101000111: data = 6'b010101;
12'b11111101001000: data = 6'b010101;
12'b11111101001001: data = 6'b010101;
12'b11111101001010: data = 6'b010101;
12'b11111101001011: data = 6'b010101;
12'b11111101001100: data = 6'b010101;
12'b11111101001101: data = 6'b010101;
12'b11111101001110: data = 6'b010101;
12'b11111101001111: data = 6'b010101;
12'b11111101010000: data = 6'b010101;
12'b11111101010001: data = 6'b010101;
12'b11111101010010: data = 6'b010101;
12'b11111101010011: data = 6'b010101;
12'b11111101010100: data = 6'b010101;
12'b11111101010101: data = 6'b010101;
12'b11111101010110: data = 6'b010101;
12'b11111101010111: data = 6'b101010;
12'b11111101011000: data = 6'b101010;
12'b11111101011001: data = 6'b101010;
12'b11111101011010: data = 6'b000000;
12'b11111101011011: data = 6'b101010;
12'b11111101011100: data = 6'b101010;
12'b11111101011101: data = 6'b101010;
12'b11111101011110: data = 6'b101010;
12'b11111101011111: data = 6'b101010;
12'b11111101100000: data = 6'b000000;
12'b11111101100001: data = 6'b000000;
12'b11111101100010: data = 6'b010101;
12'b11111101100011: data = 6'b010101;
12'b11111101100100: data = 6'b010101;
12'b11111101100101: data = 6'b010101;
12'b11111101100110: data = 6'b010101;
12'b11111101100111: data = 6'b010101;
12'b11111101101000: data = 6'b010101;
12'b11111101101001: data = 6'b010101;
12'b11111101101010: data = 6'b010101;
12'b11111101101011: data = 6'b010101;
12'b11111101101100: data = 6'b010101;
12'b11111101101101: data = 6'b010101;
12'b11111101101110: data = 6'b010101;
12'b11111101101111: data = 6'b010101;
12'b11111101110000: data = 6'b010101;
12'b11111101110001: data = 6'b010101;
12'b11111101110010: data = 6'b010101;
12'b11111101110011: data = 6'b010101;
12'b11111101110100: data = 6'b010101;
12'b11111101110101: data = 6'b010101;
12'b11111101110110: data = 6'b010101;
12'b11111101110111: data = 6'b010101;
12'b11111101111000: data = 6'b010101;
12'b11111101111001: data = 6'b010101;
12'b11111101111010: data = 6'b010101;
12'b11111101111011: data = 6'b010101;
12'b11111101111100: data = 6'b010101;
12'b11111101111101: data = 6'b010101;
12'b11111101111110: data = 6'b010101;
12'b11111101111111: data = 6'b010101;
12'b111111010000000: data = 6'b010101;
12'b111111010000001: data = 6'b010101;
12'b111111010000010: data = 6'b010101;
12'b111111010000011: data = 6'b010101;
12'b111111010000100: data = 6'b010101;
12'b111111010000101: data = 6'b101010;
12'b111111010000110: data = 6'b010101;
12'b111111010000111: data = 6'b010101;
12'b111111010001000: data = 6'b010101;
12'b111111010001001: data = 6'b101010;
12'b111111010001010: data = 6'b101010;
12'b111111010001011: data = 6'b101010;
12'b111111010001100: data = 6'b101010;
12'b111111010001101: data = 6'b010101;
12'b111111010001110: data = 6'b010101;
12'b111111010001111: data = 6'b010101;
12'b111111010010000: data = 6'b010101;
12'b111111010010001: data = 6'b010101;
12'b111111010010010: data = 6'b010101;
12'b111111010010011: data = 6'b010101;
12'b111111010010100: data = 6'b010101;
12'b111111010010101: data = 6'b010101;
12'b111111010010110: data = 6'b010101;
12'b111111010010111: data = 6'b010101;
12'b111111010011000: data = 6'b010101;
12'b111111010011001: data = 6'b010101;
12'b111111010011010: data = 6'b010101;
12'b111111010011011: data = 6'b010101;
12'b111111010011100: data = 6'b010101;
12'b111111010011101: data = 6'b010101;
12'b111111010011110: data = 6'b010101;
12'b111111010011111: data = 6'b010101;
12'b111111010100000: data = 6'b010101;
12'b111111010100001: data = 6'b010101;
12'b111111010100010: data = 6'b010101;
12'b111111010100011: data = 6'b010101;
12'b111111010100100: data = 6'b010101;
12'b111111010100101: data = 6'b010101;
12'b111111010100110: data = 6'b010101;
12'b111111010100111: data = 6'b010101;
12'b111111010101000: data = 6'b010101;
12'b111111010101001: data = 6'b010101;
12'b111111010101010: data = 6'b010101;
12'b1111111000000: data = 6'b010101;
12'b1111111000001: data = 6'b010101;
12'b1111111000010: data = 6'b010101;
12'b1111111000011: data = 6'b010101;
12'b1111111000100: data = 6'b010101;
12'b1111111000101: data = 6'b010101;
12'b1111111000110: data = 6'b010101;
12'b1111111000111: data = 6'b010101;
12'b1111111001000: data = 6'b010101;
12'b1111111001001: data = 6'b010101;
12'b1111111001010: data = 6'b010101;
12'b1111111001011: data = 6'b010101;
12'b1111111001100: data = 6'b010101;
12'b1111111001101: data = 6'b010101;
12'b1111111001110: data = 6'b010101;
12'b1111111001111: data = 6'b010101;
12'b1111111010000: data = 6'b010101;
12'b1111111010001: data = 6'b010101;
12'b1111111010010: data = 6'b010101;
12'b1111111010011: data = 6'b010101;
12'b1111111010100: data = 6'b010101;
12'b1111111010101: data = 6'b010101;
12'b1111111010110: data = 6'b010101;
12'b1111111010111: data = 6'b010101;
12'b1111111011000: data = 6'b010101;
12'b1111111011001: data = 6'b010101;
12'b1111111011010: data = 6'b010101;
12'b1111111011011: data = 6'b010101;
12'b1111111011100: data = 6'b010101;
12'b1111111011101: data = 6'b010101;
12'b1111111011110: data = 6'b010101;
12'b1111111011111: data = 6'b010101;
12'b1111111100000: data = 6'b010101;
12'b1111111100001: data = 6'b010101;
12'b1111111100010: data = 6'b010101;
12'b1111111100011: data = 6'b010101;
12'b1111111100100: data = 6'b010101;
12'b1111111100101: data = 6'b010101;
12'b1111111100110: data = 6'b010101;
12'b1111111100111: data = 6'b010101;
12'b1111111101000: data = 6'b010101;
12'b1111111101001: data = 6'b010101;
12'b1111111101010: data = 6'b010101;
12'b1111111101011: data = 6'b010101;
12'b1111111101100: data = 6'b010101;
12'b1111111101101: data = 6'b010101;
12'b1111111101110: data = 6'b010101;
12'b1111111101111: data = 6'b010101;
12'b1111111110000: data = 6'b010101;
12'b1111111110001: data = 6'b010101;
12'b1111111110010: data = 6'b010101;
12'b1111111110011: data = 6'b010101;
12'b1111111110100: data = 6'b010101;
12'b1111111110101: data = 6'b010101;
12'b1111111110110: data = 6'b010101;
12'b1111111110111: data = 6'b010101;
12'b1111111111000: data = 6'b010101;
12'b1111111111001: data = 6'b010101;
12'b1111111111010: data = 6'b010101;
12'b1111111111011: data = 6'b010101;
12'b1111111111100: data = 6'b010101;
12'b1111111111101: data = 6'b010101;
12'b1111111111110: data = 6'b010101;
12'b1111111111111: data = 6'b010101;
12'b11111111000000: data = 6'b010101;
12'b11111111000001: data = 6'b010101;
12'b11111111000010: data = 6'b010101;
12'b11111111000011: data = 6'b010101;
12'b11111111000100: data = 6'b010101;
12'b11111111000101: data = 6'b010101;
12'b11111111000110: data = 6'b010101;
12'b11111111000111: data = 6'b010101;
12'b11111111001000: data = 6'b010101;
12'b11111111001001: data = 6'b010101;
12'b11111111001010: data = 6'b010101;
12'b11111111001011: data = 6'b010101;
12'b11111111001100: data = 6'b010101;
12'b11111111001101: data = 6'b010101;
12'b11111111001110: data = 6'b010101;
12'b11111111001111: data = 6'b010101;
12'b11111111010000: data = 6'b010101;
12'b11111111010001: data = 6'b010101;
12'b11111111010010: data = 6'b010101;
12'b11111111010011: data = 6'b010101;
12'b11111111010100: data = 6'b010101;
12'b11111111010101: data = 6'b010101;
12'b11111111010110: data = 6'b010101;
12'b11111111010111: data = 6'b010101;
12'b11111111011000: data = 6'b010101;
12'b11111111011001: data = 6'b010101;
12'b11111111011010: data = 6'b010101;
12'b11111111011011: data = 6'b010101;
12'b11111111011100: data = 6'b010101;
12'b11111111011101: data = 6'b010101;
12'b11111111011110: data = 6'b010101;
12'b11111111011111: data = 6'b010101;
12'b11111111100000: data = 6'b010101;
12'b11111111100001: data = 6'b010101;
12'b11111111100010: data = 6'b010101;
12'b11111111100011: data = 6'b010101;
12'b11111111100100: data = 6'b010101;
12'b11111111100101: data = 6'b010101;
12'b11111111100110: data = 6'b010101;
12'b11111111100111: data = 6'b010101;
12'b11111111101000: data = 6'b010101;
12'b11111111101001: data = 6'b010101;
12'b11111111101010: data = 6'b010101;
12'b11111111101011: data = 6'b010101;
12'b11111111101100: data = 6'b010101;
12'b11111111101101: data = 6'b010101;
12'b11111111101110: data = 6'b010101;
12'b11111111101111: data = 6'b010101;
12'b11111111110000: data = 6'b010101;
12'b11111111110001: data = 6'b010101;
12'b11111111110010: data = 6'b010101;
12'b11111111110011: data = 6'b010101;
12'b11111111110100: data = 6'b010101;
12'b11111111110101: data = 6'b010101;
12'b11111111110110: data = 6'b010101;
12'b11111111110111: data = 6'b010101;
12'b11111111111000: data = 6'b010101;
12'b11111111111001: data = 6'b010101;
12'b11111111111010: data = 6'b010101;
12'b11111111111011: data = 6'b010101;
12'b11111111111100: data = 6'b010101;
12'b11111111111101: data = 6'b010101;
12'b11111111111110: data = 6'b010101;
12'b11111111111111: data = 6'b010101;
12'b111111110000000: data = 6'b010101;
12'b111111110000001: data = 6'b010101;
12'b111111110000010: data = 6'b010101;
12'b111111110000011: data = 6'b010101;
12'b111111110000100: data = 6'b010101;
12'b111111110000101: data = 6'b010101;
12'b111111110000110: data = 6'b010101;
12'b111111110000111: data = 6'b010101;
12'b111111110001000: data = 6'b010101;
12'b111111110001001: data = 6'b010101;
12'b111111110001010: data = 6'b010101;
12'b111111110001011: data = 6'b010101;
12'b111111110001100: data = 6'b010101;
12'b111111110001101: data = 6'b010101;
12'b111111110001110: data = 6'b010101;
12'b111111110001111: data = 6'b010101;
12'b111111110010000: data = 6'b010101;
12'b111111110010001: data = 6'b010101;
12'b111111110010010: data = 6'b010101;
12'b111111110010011: data = 6'b010101;
12'b111111110010100: data = 6'b010101;
12'b111111110010101: data = 6'b010101;
12'b111111110010110: data = 6'b010101;
12'b111111110010111: data = 6'b010101;
12'b111111110011000: data = 6'b010101;
12'b111111110011001: data = 6'b010101;
12'b111111110011010: data = 6'b010101;
12'b111111110011011: data = 6'b010101;
12'b111111110011100: data = 6'b010101;
12'b111111110011101: data = 6'b010101;
12'b111111110011110: data = 6'b010101;
12'b111111110011111: data = 6'b010101;
12'b111111110100000: data = 6'b010101;
12'b111111110100001: data = 6'b010101;
12'b111111110100010: data = 6'b010101;
12'b111111110100011: data = 6'b010101;
12'b111111110100100: data = 6'b010101;
12'b111111110100101: data = 6'b010101;
12'b111111110100110: data = 6'b010101;
12'b111111110100111: data = 6'b010101;
12'b111111110101000: data = 6'b010101;
12'b111111110101001: data = 6'b010101;
12'b111111110101010: data = 6'b010101;
    endcase
end
endmodule
